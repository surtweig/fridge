
module xcm_clk_pll (
	xcm_clk_pll_in_clk,
	xcm_clk_pll_reset_reset,
	xcm_clk_pll_out_clk);	

	input		xcm_clk_pll_in_clk;
	input		xcm_clk_pll_reset_reset;
	output		xcm_clk_pll_out_clk;
endmodule
