
module vga_pll (
	vga_pll_clk_in_clk,
	vga_pll_reset_reset,
	vga_pll_clk_out_clk);	

	input		vga_pll_clk_in_clk;
	input		vga_pll_reset_reset;
	output		vga_pll_clk_out_clk;
endmodule
