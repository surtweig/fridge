-- vga_pll.vhd

-- Generated using ACDS version 17.0 595

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity vga_pll is
	port (
		vga_pll_clk_in_clk  : in  std_logic := '0'; --  vga_pll_clk_in.clk
		vga_pll_clk_out_clk : out std_logic;        -- vga_pll_clk_out.clk
		vga_pll_reset_reset : in  std_logic := '0'  --   vga_pll_reset.reset
	);
end entity vga_pll;

architecture rtl of vga_pll is
	component vga_pll_pll_0 is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component vga_pll_pll_0;

begin

	pll_0 : component vga_pll_pll_0
		port map (
			refclk   => vga_pll_clk_in_clk,  --  refclk.clk
			rst      => vga_pll_reset_reset, --   reset.reset
			outclk_0 => vga_pll_clk_out_clk, -- outclk0.clk
			locked   => open                 -- (terminated)
		);

end architecture rtl; -- of vga_pll
