-- xcm_clk_pll.vhd

-- Generated using ACDS version 17.0 595

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity xcm_clk_pll is
	port (
		xcm_clk_pll_in_clk      : in  std_logic := '0'; --    xcm_clk_pll_in.clk
		xcm_clk_pll_out_clk     : out std_logic;        --   xcm_clk_pll_out.clk
		xcm_clk_pll_reset_reset : in  std_logic := '0'  -- xcm_clk_pll_reset.reset
	);
end entity xcm_clk_pll;

architecture rtl of xcm_clk_pll is
	component xcm_clk_pll_pll_0 is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component xcm_clk_pll_pll_0;

begin

	pll_0 : component xcm_clk_pll_pll_0
		port map (
			refclk   => xcm_clk_pll_in_clk,      --  refclk.clk
			rst      => xcm_clk_pll_reset_reset, --   reset.reset
			outclk_0 => xcm_clk_pll_out_clk,     -- outclk0.clk
			locked   => open                     -- (terminated)
		);

end architecture rtl; -- of xcm_clk_pll
