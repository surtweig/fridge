
module cpu_clk_pll (
	cpu_clk_pll_in_clk,
	cpu_clk_pll_reset_reset,
	cpu_clk_pll_out_clk);	

	input		cpu_clk_pll_in_clk;
	input		cpu_clk_pll_reset_reset;
	output		cpu_clk_pll_out_clk;
endmodule
