(
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"58", X"F0", X"43", X"F0", X"4D", X"F0", X"32", X"F0", X"20", X"F0", 
X"46", X"F0", X"72", X"F0", X"69", X"F0", X"64", X"F0", X"67", X"F0", X"65", X"F0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"20", X"B0", X"20", X"B0", 
X"20", X"B0", X"20", X"B0", X"20", X"B0", X"20", X"B0", X"2F", X"B0", X"5C", X"B0", X"20", X"B0", X"20", X"B0", 
X"20", X"B0", X"20", X"B0", X"20", X"B0", X"20", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"20", X"B0", X"5F", X"B0", 
X"5F", X"B0", X"20", X"B0", X"20", X"B0", X"20", X"B0", X"5C", X"B0", X"2F", X"B0", X"20", X"B0", X"20", X"B0", 
X"20", X"B0", X"5F", X"B0", X"5F", X"B0", X"20", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"20", X"B0", X"5C", X"B0", 
X"5F", X"B0", X"5C", X"B0", X"5F", X"B0", X"5C", X"B0", X"2F", X"B0", X"5C", X"B0", X"2F", X"B0", X"5F", X"B0", 
X"2F", X"B0", X"5F", X"B0", X"2F", X"B0", X"20", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"20", X"B0", X"20", X"B0", 
X"20", X"B0", X"5F", X"B0", X"5C", X"B0", X"5F", X"B0", X"5C", X"B0", X"2F", X"B0", X"5F", X"B0", X"2F", X"B0", 
X"5F", X"B0", X"20", X"B0", X"20", X"B0", X"20", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"20", X"B0", X"20", X"B0", 
X"5F", X"B0", X"5F", X"B0", X"2F", X"B0", X"5F", X"B0", X"2F", X"B0", X"5C", X"B0", X"5F", X"B0", X"5C", X"B0", 
X"5F", X"B0", X"5F", X"B0", X"20", X"B0", X"20", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"20", X"B0", X"2F", X"B0", 
X"5F", X"B0", X"2F", X"B0", X"20", X"B0", X"2F", X"B0", X"5C", X"B0", X"2F", X"B0", X"5C", X"B0", X"20", X"B0", 
X"5C", X"B0", X"5F", X"B0", X"5C", X"B0", X"20", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"20", X"B0", X"20", X"B0", 
X"20", X"B0", X"20", X"B0", X"20", X"B0", X"20", X"B0", X"2F", X"B0", X"5C", X"B0", X"20", X"B0", X"20", X"B0", 
X"20", X"B0", X"20", X"B0", X"20", X"B0", X"20", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"20", X"B0", X"20", X"B0", 
X"20", X"B0", X"20", X"B0", X"20", X"B0", X"20", X"B0", X"5C", X"B0", X"2F", X"B0", X"20", X"B0", X"20", X"B0", 
X"20", X"B0", X"20", X"B0", X"20", X"B0", X"20", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"50", X"F0", X"6C", X"F0", X"75", X"F0", 
X"73", X"F0", X"26", X"F0", X"4D", X"F0", X"69", X"F0", X"6E", X"F0", X"75", X"F0", X"73", X"F0", X"20", X"F0", 
X"49", X"F0", X"6E", X"F0", X"63", X"F0", X"2E", X"F0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", X"00", X"B0", 
others => 0);