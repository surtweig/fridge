library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.FridgeGlobals.all;

package FridgeWelcomeScreen is

constant WelcomeScreenData : XCM2_RAM:= 
(
X"46", X"27", X"72", X"38", X"69", X"49", X"64", X"5A", X"67", X"6B", X"65", X"7C", X"20", X"8D", X"69", X"9E", 
X"73", X"AF", X"20", X"B0", X"61", X"C1", X"20", X"D2", X"38", X"E3", X"2D", X"F4", X"62", X"05", X"69", X"16", 
X"74", X"27", X"20", X"38", X"63", X"49", X"6F", X"5A", X"6D", X"6B", X"70", X"7C", X"75", X"8D", X"74", X"9E", 
X"65", X"AF", X"72", X"B0", X"20", X"C1", X"62", X"D2", X"61", X"E3", X"73", X"F4", X"65", X"05", X"64", X"16", 
X"20", X"27", X"6F", X"38", X"6E", X"49", X"20", X"5A", X"65", X"6B", X"78", X"7C", X"74", X"8D", X"65", X"9E", 
X"6E", X"AF", X"64", X"B0", X"65", X"C1", X"64", X"D2", X"20", X"E3", X"49", X"F4", X"6E", X"05", X"74", X"16", 
X"65", X"27", X"6C", X"38", X"20", X"49", X"38", X"5A", X"30", X"6B", X"38", X"7C", X"30", X"8D", X"20", X"9E", 
X"69", X"AF", X"6E", X"B0", X"73", X"C1", X"74", X"D2", X"72", X"E3", X"75", X"F4", X"63", X"05", X"74", X"16", 
X"69", X"27", X"6F", X"38", X"6E", X"49", X"20", X"5A", X"73", X"6B", X"65", X"7C", X"74", X"8D", X"20", X"9E", 
X"77", X"AF", X"69", X"B0", X"74", X"C1", X"68", X"D2", X"20", X"E3", X"67", X"F4", X"72", X"05", X"61", X"16", 
X"70", X"27", X"68", X"38", X"69", X"49", X"63", X"5A", X"73", X"6B", X"20", X"7C", X"61", X"8D", X"63", X"9E", 
X"63", X"AF", X"65", X"B0", X"6C", X"C1", X"65", X"D2", X"72", X"E3", X"61", X"F4", X"74", X"05", X"69", X"16", 
X"6F", X"27", X"6E", X"38", X"2E", X"49", X"20", X"5A", X"43", X"6B", X"75", X"7C", X"72", X"8D", X"72", X"9E", 
X"65", X"AF", X"6E", X"B0", X"74", X"C1", X"20", X"D2", X"69", X"E3", X"6D", X"F4", X"70", X"05", X"6C", X"16", 
X"65", X"27", X"6D", X"38", X"65", X"49", X"6E", X"5A", X"74", X"6B", X"61", X"7C", X"74", X"8D", X"69", X"9E", 
X"6F", X"AF", X"6E", X"B0", X"20", X"C1", X"63", X"D2", X"6F", X"E3", X"6E", X"F4", X"73", X"05", X"69", X"16", 
X"73", X"27", X"74", X"38", X"73", X"49", X"20", X"5A", X"6F", X"6B", X"66", X"7C", X"20", X"8D", X"61", X"9E", 
X"6E", X"AF", X"20", X"B0", X"65", X"C1", X"6D", X"D2", X"75", X"E3", X"6C", X"F4", X"61", X"05", X"74", X"16", 
X"6F", X"27", X"72", X"38", X"20", X"49", X"28", X"5A", X"57", X"6B", X"69", X"7C", X"6E", X"8D", X"64", X"9E", 
X"6F", X"AF", X"77", X"B0", X"73", X"C1", X"20", X"D2", X"78", X"E3", X"36", X"F4", X"34", X"05", X"20", X"16", 
X"2B", X"27", X"20", X"38", X"44", X"49", X"69", X"5A", X"72", X"6B", X"65", X"7C", X"63", X"8D", X"74", X"9E", 
X"58", X"AF", X"20", X"B0", X"31", X"C1", X"31", X"D2", X"29", X"E3", X"20", X"F4", X"61", X"05", X"6E", X"16", 
X"64", X"27", X"20", X"38", X"56", X"49", X"48", X"5A", X"44", X"6B", X"4C", X"7C", X"20", X"8D", X"64", X"9E", 
X"65", X"AF", X"73", X"B0", X"69", X"C1", X"67", X"D2", X"6E", X"E3", X"20", X"F4", X"66", X"05", X"6F", X"16", 
X"72", X"27", X"20", X"38", X"46", X"49", X"50", X"5A", X"47", X"6B", X"41", X"7C", X"20", X"8D", X"64", X"9E", 
X"65", X"AF", X"76", X"B0", X"65", X"C1", X"6C", X"D2", X"6F", X"E3", X"70", X"F4", X"6D", X"05", X"65", X"16", 
X"6E", X"27", X"74", X"38", X"20", X"49", X"62", X"5A", X"6F", X"6B", X"61", X"7C", X"72", X"8D", X"64", X"9E", 
X"20", X"AF", X"54", X"B0", X"65", X"C1", X"72", X"D2", X"61", X"E3", X"73", X"F4", X"69", X"05", X"63", X"16", 
X"20", X"27", X"44", X"38", X"45", X"49", X"30", X"5A", X"2D", X"6B", X"43", X"7C", X"56", X"8D", X"20", X"9E", 
X"28", X"AF", X"41", X"B0", X"6C", X"C1", X"74", X"D2", X"65", X"E3", X"72", X"F4", X"61", X"05", X"20", X"16", 
X"43", X"27", X"79", X"38", X"63", X"49", X"6C", X"5A", X"6F", X"6B", X"6E", X"7C", X"65", X"8D", X"20", X"9E", 
X"56", X"AF", X"29", X"B0", X"2C", X"C1", X"20", X"D2", X"61", X"E3", X"73", X"F4", X"20", X"05", X"77", X"16", 
X"65", X"27", X"6C", X"38", X"6C", X"49", X"20", X"5A", X"61", X"6B", X"73", X"7C", X"20", X"8D", X"76", X"9E", 
X"61", X"AF", X"72", X"B0", X"69", X"C1", X"6F", X"D2", X"75", X"E3", X"73", X"F4", X"20", X"05", X"74", X"16", 
X"6F", X"27", X"6F", X"38", X"6C", X"49", X"73", X"5A", X"20", X"6B", X"73", X"7C", X"75", X"8D", X"63", X"9E", 
X"68", X"AF", X"20", X"B0", X"61", X"C1", X"73", X"D2", X"20", X"E3", X"2D", X"F4", X"20", X"05", X"61", X"16", 
X"73", X"27", X"73", X"38", X"65", X"49", X"6D", X"5A", X"62", X"6B", X"6C", X"7C", X"79", X"8D", X"20", X"9E", 
X"63", X"AF", X"6F", X"B0", X"6D", X"C1", X"70", X"D2", X"69", X"E3", X"6C", X"F4", X"65", X"05", X"72", X"16", 
X"2C", X"27", X"20", X"38", X"63", X"49", X"75", X"5A", X"73", X"6B", X"74", X"7C", X"6F", X"8D", X"6D", X"9E", 
X"20", X"AF", X"73", X"B0", X"69", X"C1", X"6D", X"D2", X"70", X"E3", X"6C", X"F4", X"69", X"05", X"73", X"16", 
X"74", X"27", X"69", X"38", X"63", X"49", X"20", X"5A", X"6C", X"6B", X"61", X"7C", X"6E", X"8D", X"67", X"9E", 
X"75", X"AF", X"61", X"B0", X"67", X"C1", X"65", X"D2", X"20", X"E3", X"63", X"F4", X"6F", X"05", X"6D", X"16", 
X"70", X"27", X"69", X"38", X"6C", X"49", X"65", X"5A", X"72", X"6B", X"20", X"7C", X"61", X"8D", X"6E", X"9E", 
X"64", X"AF", X"20", X"B0", X"61", X"C1", X"6E", X"D2", X"20", X"E3", X"49", X"F4", X"44", X"05", X"45", X"16", 
X"2E", X"27", X"53", X"38", X"79", X"49", X"73", X"5A", X"74", X"6B", X"65", X"7C", X"6D", X"8D", X"20", X"9E", 
X"73", X"AF", X"70", X"B0", X"65", X"C1", X"63", X"D2", X"73", X"E3", X"20", X"F4", X"43", X"05", X"50", X"16", 
X"55", X"27", X"20", X"38", X"4D", X"49", X"6F", X"5A", X"64", X"6B", X"69", X"7C", X"66", X"8D", X"69", X"9E", 
X"65", X"AF", X"64", X"B0", X"20", X"C1", X"42", X"D2", X"69", X"E3", X"67", X"F4", X"2D", X"05", X"45", X"16", 
X"6E", X"27", X"64", X"38", X"69", X"49", X"61", X"5A", X"6E", X"6B", X"20", X"7C", X"49", X"8D", X"6E", X"9E", 
X"74", X"AF", X"65", X"B0", X"6C", X"C1", X"20", X"D2", X"38", X"E3", X"30", X"F4", X"38", X"05", X"30", X"16", 
X"20", X"27", X"47", X"38", X"72", X"49", X"61", X"5A", X"70", X"6B", X"68", X"7C", X"69", X"8D", X"63", X"9E", 
X"61", X"AF", X"6C", X"B0", X"20", X"C1", X"69", X"D2", X"6E", X"E3", X"73", X"F4", X"74", X"05", X"72", X"16", 
X"75", X"27", X"63", X"38", X"74", X"49", X"69", X"5A", X"6F", X"6B", X"6E", X"7C", X"73", X"8D", X"20", X"9E", 
X"31", X"AF", X"30", X"B0", X"20", X"C1", X"4D", X"D2", X"48", X"E3", X"7A", X"F4", X"20", X"05", X"63", X"16", 
X"6C", X"27", X"6F", X"38", X"63", X"49", X"6B", X"5A", X"20", X"6B", X"66", X"7C", X"72", X"8D", X"65", X"9E", 
X"71", X"AF", X"75", X"B0", X"65", X"C1", X"6E", X"D2", X"63", X"E3", X"79", X"F4", X"20", X"05", X"52", X"16", 
X"41", X"27", X"4D", X"38", X"20", X"49", X"36", X"5A", X"34", X"6B", X"20", X"7C", X"4B", X"8D", X"42", X"9E", 
X"20", X"AF", X"28", X"B0", X"31", X"C1", X"36", X"D2", X"2D", X"E3", X"62", X"F4", X"69", X"05", X"74", X"16", 
X"20", X"27", X"61", X"38", X"64", X"49", X"64", X"5A", X"72", X"6B", X"65", X"7C", X"73", X"8D", X"73", X"9E", 
X"29", X"AF", X"20", X"B0", X"56", X"C1", X"69", X"D2", X"64", X"E3", X"65", X"F4", X"6F", X"05", X"20", X"16", 
X"44", X"27", X"69", X"38", X"73", X"49", X"70", X"5A", X"6C", X"6B", X"61", X"7C", X"79", X"8D", X"3A", X"9E", 
X"20", X"AF", X"32", X"B0", X"34", X"C1", X"30", X"D2", X"78", X"E3", X"31", X"F4", X"36", X"05", X"30", X"16", 
X"20", X"27", X"70", X"38", X"69", X"49", X"78", X"5A", X"65", X"6B", X"6C", X"7C", X"73", X"8D", X"20", X"9E", 
X"34", X"AF", X"2D", X"B0", X"62", X"C1", X"69", X"D2", X"74", X"E3", X"20", X"F4", X"70", X"05", X"61", X"16", 
X"6C", X"27", X"6C", X"38", X"65", X"49", X"74", X"5A", X"74", X"6B", X"65", X"7C", X"20", X"8D", X"28", X"9E", 
X"31", X"AF", X"36", X"B0", X"20", X"C1", X"63", X"D2", X"6F", X"E3", X"6C", X"F4", X"6F", X"05", X"72", X"16", 
X"73", X"27", X"29", X"38", X"20", X"49", X"66", X"5A", X"72", X"6B", X"6F", X"7C", X"6D", X"8D", X"20", X"9E", 
X"34", X"AF", X"30", X"B0", X"39", X"C1", X"36", X"D2", X"20", X"E3", X"70", X"F4", X"6F", X"05", X"73", X"16", 
X"73", X"27", X"69", X"38", X"62", X"49", X"6C", X"5A", X"65", X"6B", X"20", X"7C", X"63", X"8D", X"6F", X"9E", 
X"6C", X"AF", X"6F", X"B0", X"72", X"C1", X"73", X"D2", X"20", X"E3", X"54", X"F4", X"77", X"05", X"6F", X"16", 
X"20", X"27", X"66", X"38", X"72", X"49", X"61", X"5A", X"6D", X"6B", X"65", X"7C", X"62", X"8D", X"75", X"9E", 
X"66", X"AF", X"66", X"B0", X"65", X"C1", X"72", X"D2", X"73", X"E3", X"20", X"F4", X"32", X"05", X"34", X"16", 
X"30", X"27", X"78", X"38", X"31", X"49", X"36", X"5A", X"30", X"6B", X"78", X"7C", X"34", X"8D", X"20", X"9E", 
X"36", X"AF", X"34", X"B0", X"20", X"C1", X"4B", X"D2", X"42", X"E3", X"20", X"F4", X"73", X"05", X"70", X"16", 
X"72", X"27", X"69", X"38", X"74", X"49", X"65", X"5A", X"20", X"6B", X"6D", X"7C", X"65", X"8D", X"6D", X"9E", 
X"6F", X"AF", X"72", X"B0", X"79", X"C1", X"20", X"D2", X"28", X"E3", X"31", X"F4", X"30", X"05", X"32", X"16", 
X"20", X"27", X"4B", X"38", X"42", X"49", X"20", X"5A", X"74", X"6B", X"6F", X"7C", X"74", X"8D", X"61", X"9E", 
X"6C", X"AF", X"20", X"B0", X"76", X"C1", X"69", X"D2", X"64", X"E3", X"65", X"F4", X"6F", X"05", X"20", X"16", 
X"6D", X"27", X"65", X"38", X"6D", X"49", X"6F", X"5A", X"72", X"6B", X"79", X"7C", X"29", X"8D", X"20", X"9E", 
X"34", X"AF", X"30", X"B0", X"78", X"C1", X"32", X"D2", X"30", X"E3", X"20", X"F4", X"41", X"05", X"53", X"16", 
X"43", X"27", X"49", X"38", X"49", X"49", X"20", X"5A", X"74", X"6B", X"65", X"7C", X"78", X"8D", X"74", X"9E", 
X"20", X"AF", X"6D", X"B0", X"6F", X"C1", X"64", X"D2", X"65", X"E3", X"20", X"F4", X"28", X"05", X"36", X"16", 
X"78", X"27", X"38", X"38", X"20", X"49", X"66", X"5A", X"6F", X"6B", X"6E", X"7C", X"74", X"8D", X"29", X"9E", 
X"20", X"AF", X"52", X"B0", X"4F", X"C1", X"4D", X"D2", X"20", X"E3", X"53", X"F4", X"44", X"05", X"20", X"16", 
X"63", X"27", X"61", X"38", X"72", X"49", X"64", X"5A", X"20", X"6B", X"28", X"7C", X"31", X"8D", X"36", X"9E", 
X"20", X"AF", X"4D", X"B0", X"42", X"C1", X"20", X"D2", X"6D", X"E3", X"61", X"F4", X"78", X"05", X"69", X"16", 
X"6D", X"27", X"75", X"38", X"6D", X"49", X"29", X"5A", X"80", X"80", X"80", X"80", X"80", X"88", X"47", X"47", 
X"77", X"47", X"47", X"67", X"67", X"88", X"48", X"05", X"84", X"86", X"64", X"74", X"76", X"76", X"57", X"88", 
X"00", X"87", X"7F", X"93", X"93", X"83", X"83", X"88", X"09", X"00", X"09", X"00", X"00", X"90", X"00", X"80", 
X"30", X"80", X"80", X"90", X"00", X"80", X"90", X"00", X"18", X"03", X"08", X"00", X"03", X"08", X"08", X"08", 
X"77", X"77", X"77", X"77", X"87", X"77", X"27", X"87", X"78", X"02", X"77", X"87", X"77", X"77", X"77", X"87", 
X"78", X"77", X"77", X"77", X"77", X"87", X"78", X"77", X"87", X"27", X"77", X"77", X"72", X"88", X"77", X"87", 
X"77", X"78", X"77", X"88", X"88", X"88", X"08", X"06", X"00", X"08", X"00", X"80", X"00", X"00", X"00", X"08", 
X"08", X"00", X"00", X"02", X"08", X"88", X"20", X"88", X"00", X"00", X"00", X"00", X"88", X"48", X"80", X"80", 
X"80", X"50", X"84", X"05", X"08", X"04", X"74", X"7C", X"47", X"47", X"56", X"74", X"74", X"70", X"00", X"08", 
X"85", X"84", X"77", X"47", X"56", X"78", X"78", X"80", X"50", X"89", X"3F", X"77", X"78", X"38", X"98", X"90", 
X"80", X"88", X"00", X"09", X"00", X"00", X"88", X"09", X"00", X"80", X"80", X"00", X"80", X"00", X"00", X"80", 
X"80", X"10", X"09", X"08", X"00", X"08", X"00", X"00", X"77", X"78", X"77", X"77", X"77", X"77", X"77", X"27", 
X"80", X"00", X"67", X"87", X"87", X"87", X"77", X"87", X"77", X"78", X"77", X"77", X"77", X"77", X"77", X"77", 
X"77", X"77", X"77", X"77", X"77", X"28", X"78", X"87", X"88", X"77", X"87", X"87", X"70", X"20", X"68", X"08", 
X"08", X"08", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"80", X"00", X"00", X"00", X"00", X"02", X"08", 
X"08", X"00", X"00", X"10", X"08", X"08", X"80", X"84", X"08", X"08", X"08", X"00", X"48", X"85", X"74", X"77", 
X"74", X"74", X"74", X"74", X"75", X"80", X"00", X"00", X"04", X"84", X"74", X"76", X"76", X"58", X"85", X"80", 
X"00", X"08", X"38", X"38", X"88", X"83", X"03", X"88", X"03", X"18", X"80", X"08", X"08", X"00", X"00", X"00", 
X"00", X"90", X"00", X"00", X"08", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"08", X"00", 
X"77", X"77", X"78", X"77", X"27", X"77", X"78", X"77", X"80", X"88", X"08", X"08", X"77", X"77", X"77", X"77", 
X"87", X"87", X"77", X"77", X"77", X"77", X"77", X"72", X"78", X"77", X"87", X"78", X"78", X"80", X"20", X"08", 
X"87", X"77", X"72", X"88", X"68", X"60", X"80", X"80", X"80", X"80", X"00", X"00", X"08", X"00", X"80", X"80", 
X"08", X"00", X"00", X"00", X"00", X"08", X"00", X"83", X"08", X"08", X"00", X"08", X"88", X"80", X"48", X"08", 
X"08", X"08", X"08", X"08", X"00", X"47", X"47", X"C7", X"44", X"74", X"7C", X"77", X"47", X"40", X"00", X"00", 
X"00", X"45", X"67", X"C7", X"57", X"78", X"80", X"08", X"08", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
X"00", X"00", X"00", X"00", X"00", X"08", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"80", X"00", 
X"00", X"00", X"00", X"00", X"80", X"00", X"00", X"00", X"87", X"77", X"77", X"77", X"77", X"77", X"78", X"77", 
X"80", X"80", X"80", X"80", X"77", X"87", X"87", X"87", X"77", X"78", X"77", X"77", X"87", X"87", X"77", X"77", 
X"28", X"88", X"87", X"72", X"78", X"88", X"88", X"88", X"87", X"77", X"78", X"82", X"80", X"80", X"60", X"80", 
X"80", X"80", X"00", X"00", X"00", X"00", X"00", X"08", X"00", X"08", X"00", X"00", X"00", X"00", X"00", X"03", 
X"03", X"01", X"80", X"00", X"80", X"80", X"80", X"88", X"04", X"08", X"08", X"05", X"08", X"74", X"74", X"74", 
X"74", X"74", X"74", X"74", X"75", X"00", X"00", X"00", X"07", X"67", X"47", X"47", X"48", X"48", X"80", X"00", 
X"50", X"80", X"00", X"80", X"10", X"08", X"00", X"08", X"00", X"00", X"08", X"08", X"01", X"00", X"08", X"08", 
X"00", X"00", X"80", X"80", X"08", X"00", X"01", X"80", X"80", X"80", X"08", X"00", X"00", X"90", X"08", X"00", 
X"77", X"78", X"77", X"77", X"78", X"78", X"77", X"67", X"72", X"06", X"08", X"08", X"77", X"77", X"77", X"78", 
X"78", X"27", X"77", X"87", X"87", X"77", X"77", X"77", X"77", X"27", X"88", X"88", X"88", X"28", X"88", X"08", 
X"87", X"78", X"88", X"88", X"68", X"68", X"08", X"88", X"80", X"08", X"06", X"86", X"06", X"06", X"06", X"06", 
X"08", X"00", X"00", X"00", X"80", X"00", X"80", X"00", X"00", X"00", X"00", X"00", X"88", X"88", X"88", X"50", 
X"80", X"80", X"84", X"08", X"08", X"87", X"47", X"47", X"47", X"45", X"67", X"56", X"78", X"00", X"00", X"00", 
X"45", X"67", X"47", X"47", X"87", X"50", X"00", X"00", X"00", X"00", X"80", X"00", X"80", X"00", X"01", X"00", 
X"08", X"08", X"00", X"00", X"00", X"80", X"00", X"00", X"08", X"00", X"01", X"00", X"00", X"10", X"00", X"00", 
X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"77", X"77", X"87", X"87", X"77", X"77", X"77", X"78", 
X"78", X"88", X"88", X"08", X"88", X"77", X"87", X"78", X"77", X"78", X"77", X"77", X"87", X"28", X"78", X"77", 
X"78", X"88", X"28", X"88", X"88", X"88", X"82", X"80", X"87", X"88", X"78", X"88", X"80", X"88", X"08", X"88", 
X"88", X"80", X"60", X"60", X"68", X"60", X"68", X"00", X"60", X"68", X"08", X"00", X"00", X"80", X"08", X"08", 
X"00", X"00", X"90", X"00", X"50", X"80", X"80", X"80", X"80", X"58", X"08", X"08", X"08", X"47", X"47", X"C7", 
X"47", X"47", X"47", X"65", X"65", X"00", X"05", X"08", X"47", X"46", X"57", X"65", X"88", X"80", X"58", X"00", 
X"00", X"01", X"08", X"00", X"80", X"08", X"00", X"80", X"01", X"00", X"01", X"08", X"00", X"08", X"00", X"80", 
X"00", X"80", X"00", X"08", X"00", X"80", X"08", X"00", X"10", X"08", X"01", X"08", X"00", X"08", X"00", X"80", 
X"77", X"77", X"77", X"78", X"77", X"27", X"78", X"88", X"88", X"08", X"02", X"08", X"08", X"77", X"77", X"80", 
X"88", X"77", X"78", X"72", X"78", X"77", X"72", X"77", X"20", X"88", X"00", X"60", X"28", X"88", X"88", X"08", 
X"08", X"83", X"88", X"68", X"86", X"80", X"87", X"88", X"88", X"84", X"86", X"66", X"86", X"86", X"06", X"68", 
X"00", X"00", X"00", X"00", X"00", X"02", X"00", X"00", X"09", X"00", X"00", X"00", X"80", X"88", X"08", X"88", 
X"08", X"00", X"80", X"80", X"48", X"84", X"74", X"74", X"74", X"84", X"74", X"78", X"80", X"00", X"00", X"04", 
X"74", X"74", X"74", X"78", X"48", X"00", X"00", X"08", X"00", X"00", X"00", X"00", X"00", X"00", X"08", X"00", 
X"00", X"08", X"00", X"00", X"01", X"00", X"10", X"00", X"80", X"00", X"80", X"00", X"00", X"00", X"00", X"08", 
X"00", X"00", X"00", X"00", X"08", X"00", X"00", X"00", X"87", X"77", X"72", X"78", X"77", X"87", X"78", X"00", 
X"02", X"88", X"80", X"88", X"88", X"88", X"77", X"20", X"60", X"87", X"77", X"78", X"78", X"87", X"77", X"87", 
X"72", X"02", X"00", X"88", X"06", X"82", X"02", X"02", X"83", X"68", X"78", X"88", X"88", X"88", X"88", X"78", 
X"88", X"84", X"86", X"86", X"66", X"66", X"06", X"66", X"66", X"66", X"68", X"08", X"00", X"00", X"80", X"80", 
X"00", X"00", X"01", X"00", X"88", X"04", X"80", X"04", X"08", X"08", X"08", X"08", X"08", X"84", X"74", X"74", 
X"86", X"54", X"76", X"54", X"80", X"80", X"00", X"74", X"74", X"74", X"84", X"88", X"80", X"00", X"00", X"00", 
X"80", X"80", X"08", X"00", X"80", X"80", X"00", X"00", X"80", X"00", X"00", X"80", X"00", X"80", X"00", X"00", 
X"08", X"00", X"00", X"08", X"00", X"80", X"80", X"00", X"08", X"00", X"80", X"80", X"00", X"08", X"08", X"00", 
X"77", X"77", X"77", X"72", X"78", X"88", X"80", X"88", X"88", X"06", X"88", X"82", X"88", X"80", X"88", X"08", 
X"80", X"87", X"77", X"77", X"77", X"27", X"87", X"27", X"80", X"88", X"02", X"68", X"88", X"86", X"08", X"60", 
X"88", X"87", X"87", X"78", X"88", X"87", X"78", X"87", X"88", X"46", X"46", X"68", X"48", X"66", X"66", X"86", 
X"68", X"60", X"86", X"00", X"00", X"00", X"00", X"00", X"00", X"80", X"80", X"01", X"88", X"80", X"08", X"80", 
X"80", X"40", X"85", X"08", X"05", X"67", X"47", X"47", X"47", X"47", X"47", X"48", X"00", X"00", X"05", X"47", 
X"47", X"47", X"48", X"85", X"00", X"08", X"00", X"50", X"00", X"00", X"80", X"00", X"10", X"00", X"80", X"80", 
X"00", X"18", X"00", X"00", X"80", X"00", X"80", X"80", X"00", X"08", X"01", X"00", X"00", X"00", X"00", X"80", 
X"00", X"00", X"00", X"00", X"10", X"00", X"00", X"08", X"77", X"78", X"77", X"78", X"78", X"20", X"86", X"08", 
X"88", X"88", X"86", X"88", X"68", X"86", X"86", X"88", X"60", X"87", X"87", X"77", X"77", X"77", X"78", X"02", 
X"80", X"28", X"00", X"02", X"88", X"88", X"02", X"06", X"88", X"77", X"87", X"88", X"88", X"87", X"77", X"88", 
X"88", X"88", X"48", X"46", X"66", X"66", X"86", X"68", X"66", X"66", X"66", X"66", X"80", X"00", X"00", X"08", 
X"00", X"90", X"00", X"00", X"80", X"80", X"80", X"80", X"80", X"80", X"08", X"08", X"08", X"84", X"76", X"54", 
X"84", X"74", X"74", X"88", X"00", X"80", X"04", X"76", X"56", X"58", X"48", X"80", X"80", X"00", X"00", X"00", 
X"05", X"00", X"08", X"00", X"08", X"00", X"01", X"00", X"80", X"00", X"81", X"00", X"08", X"00", X"10", X"00", 
X"00", X"00", X"00", X"80", X"80", X"08", X"00", X"10", X"80", X"18", X"00", X"80", X"08", X"00", X"80", X"00", 
X"78", X"77", X"88", X"80", X"68", X"88", X"08", X"88", X"77", X"77", X"77", X"88", X"76", X"88", X"88", X"88", 
X"08", X"08", X"77", X"87", X"77", X"78", X"88", X"00", X"06", X"02", X"08", X"88", X"88", X"20", X"00", X"02", 
X"87", X"77", X"77", X"88", X"08", X"77", X"87", X"88", X"84", X"66", X"66", X"74", X"74", X"74", X"66", X"74", 
X"67", X"68", X"68", X"68", X"60", X"00", X"00", X"00", X"80", X"00", X"90", X"00", X"88", X"05", X"08", X"08", 
X"08", X"08", X"04", X"08", X"08", X"47", X"47", X"68", X"47", X"47", X"47", X"48", X"00", X"00", X"88", X"47", 
X"68", X"68", X"80", X"00", X"00", X"80", X"80", X"80", X"00", X"00", X"00", X"08", X"00", X"10", X"00", X"00", 
X"00", X"80", X"00", X"00", X"00", X"08", X"00", X"80", X"80", X"08", X"00", X"00", X"00", X"10", X"00", X"00", 
X"00", X"00", X"00", X"00", X"00", X"01", X"00", X"00", X"77", X"28", X"02", X"88", X"88", X"82", X"86", X"87", 
X"77", X"77", X"77", X"78", X"88", X"68", X"68", X"68", X"68", X"60", X"87", X"87", X"87", X"77", X"28", X"80", 
X"20", X"86", X"87", X"67", X"60", X"80", X"68", X"08", X"87", X"77", X"57", X"88", X"88", X"77", X"87", X"88", 
X"88", X"74", X"76", X"47", X"64", X"76", X"74", X"67", X"66", X"66", X"68", X"66", X"86", X"88", X"00", X"00", 
X"00", X"00", X"00", X"10", X"08", X"88", X"04", X"05", X"80", X"80", X"80", X"80", X"88", X"57", X"C7", X"48", 
X"65", X"74", X"74", X"80", X"00", X"00", X"8C", X"74", X"74", X"84", X"08", X"00", X"00", X"00", X"00", X"00", 
X"80", X"80", X"80", X"00", X"00", X"80", X"08", X"08", X"00", X"08", X"00", X"80", X"80", X"00", X"00", X"00", 
X"10", X"00", X"08", X"00", X"80", X"00", X"80", X"80", X"08", X"00", X"80", X"08", X"08", X"00", X"08", X"00", 
X"77", X"77", X"88", X"67", X"76", X"88", X"88", X"86", X"88", X"77", X"87", X"87", X"68", X"87", X"87", X"78", 
X"28", X"82", X"06", X"02", X"77", X"77", X"80", X"20", X"00", X"82", X"87", X"78", X"02", X"02", X"00", X"88", 
X"77", X"77", X"77", X"80", X"88", X"75", X"78", X"88", X"46", X"47", X"46", X"74", X"67", X"C6", X"7C", X"74", 
X"74", X"74", X"74", X"68", X"48", X"60", X"00", X"00", X"80", X"00", X"80", X"00", X"88", X"40", X"88", X"08", 
X"04", X"08", X"08", X"04", X"04", X"74", X"74", X"74", X"84", X"74", X"57", X"40", X"80", X"00", X"57", X"47", 
X"58", X"80", X"00", X"05", X"00", X"80", X"08", X"00", X"00", X"10", X"00", X"10", X"00", X"00", X"00", X"00", 
X"00", X"00", X"00", X"00", X"00", X"80", X"00", X"00", X"08", X"00", X"00", X"10", X"00", X"80", X"00", X"00", 
X"00", X"00", X"00", X"00", X"00", X"08", X"00", X"00", X"78", X"88", X"87", X"77", X"77", X"78", X"68", X"88", 
X"88", X"68", X"67", X"87", X"82", X"86", X"86", X"76", X"78", X"68", X"88", X"08", X"88", X"72", X"80", X"80", 
X"20", X"08", X"88", X"28", X"06", X"08", X"08", X"87", X"75", X"77", X"77", X"80", X"87", X"78", X"88", X"48", 
X"88", X"64", X"76", X"C7", X"66", X"76", X"67", X"64", X"74", X"76", X"47", X"66", X"48", X"68", X"00", X"00", 
X"08", X"00", X"10", X"80", X"08", X"88", X"08", X"08", X"08", X"08", X"08", X"08", X"88", X"47", X"76", X"54", 
X"74", X"76", X"65", X"80", X"00", X"80", X"87", X"67", X"40", X"50", X"80", X"00", X"00", X"00", X"10", X"08", 
X"00", X"08", X"00", X"08", X"08", X"00", X"80", X"01", X"80", X"08", X"00", X"50", X"01", X"00", X"80", X"80", 
X"00", X"08", X"00", X"00", X"00", X"00", X"00", X"80", X"80", X"08", X"01", X"80", X"00", X"00", X"08", X"00", 
X"80", X"28", X"77", X"77", X"76", X"77", X"88", X"68", X"60", X"88", X"77", X"77", X"87", X"87", X"88", X"68", 
X"86", X"88", X"68", X"02", X"08", X"77", X"72", X"08", X"00", X"62", X"06", X"86", X"20", X"02", X"06", X"87", 
X"87", X"87", X"58", X"80", X"88", X"87", X"88", X"06", X"46", X"74", X"67", X"64", X"7C", X"7C", X"7C", X"76", 
X"7C", X"67", X"64", X"76", X"84", X"68", X"80", X"00", X"00", X"80", X"00", X"10", X"88", X"88", X"88", X"88", 
X"08", X"05", X"08", X"00", X"85", X"67", X"C7", X"48", X"48", X"45", X"76", X"80", X"50", X"00", X"84", X"58", 
X"80", X"00", X"00", X"80", X"80", X"00", X"08", X"00", X"00", X"00", X"08", X"00", X"00", X"00", X"00", X"00", 
X"00", X"80", X"00", X"00", X"00", X"00", X"00", X"00", X"80", X"00", X"08", X"08", X"00", X"80", X"00", X"01", 
X"00", X"00", X"00", X"00", X"80", X"00", X"00", X"08", X"88", X"77", X"77", X"F7", X"77", X"77", X"78", X"88", 
X"86", X"88", X"67", X"78", X"78", X"68", X"67", X"86", X"86", X"76", X"86", X"80", X"60", X"26", X"78", X"60", 
X"20", X"02", X"88", X"80", X"28", X"02", X"08", X"87", X"88", X"77", X"78", X"88", X"78", X"88", X"88", X"88", 
X"76", X"47", X"47", X"C7", X"67", X"67", X"67", X"C7", X"67", X"47", X"47", X"46", X"84", X"84", X"60", X"00", 
X"00", X"80", X"80", X"00", X"08", X"04", X"80", X"84", X"08", X"08", X"08", X"80", X"88", X"47", X"47", X"48", 
X"57", X"66", X"54", X"00", X"00", X"00", X"00", X"88", X"08", X"00", X"00", X"00", X"00", X"80", X"00", X"00", 
X"80", X"80", X"00", X"08", X"00", X"80", X"80", X"08", X"00", X"00", X"08", X"00", X"80", X"80", X"10", X"00", 
X"01", X"80", X"00", X"00", X"00", X"01", X"80", X"00", X"08", X"00", X"80", X"00", X"01", X"08", X"00", X"00", 
X"87", X"7F", X"7F", X"67", X"F7", X"76", X"77", X"68", X"88", X"86", X"87", X"77", X"68", X"88", X"68", X"68", 
X"88", X"68", X"26", X"88", X"08", X"00", X"28", X"78", X"08", X"08", X"02", X"08", X"00", X"80", X"86", X"78", 
X"88", X"87", X"88", X"08", X"88", X"88", X"04", X"04", X"66", X"74", X"66", X"7C", X"7C", X"67", X"C7", X"66", 
X"7C", X"76", X"74", X"74", X"67", X"48", X"80", X"00", X"00", X"00", X"00", X"90", X"88", X"88", X"88", X"08", 
X"80", X"40", X"80", X"40", X"85", X"67", X"47", X"40", X"46", X"56", X"74", X"80", X"08", X"00", X"80", X"00", 
X"00", X"05", X"00", X"80", X"08", X"00", X"80", X"80", X"00", X"00", X"80", X"01", X"00", X"00", X"00", X"00", 
X"50", X"08", X"00", X"00", X"00", X"00", X"80", X"00", X"00", X"00", X"08", X"01", X"08", X"00", X"00", X"80", 
X"00", X"00", X"00", X"10", X"80", X"00", X"08", X"00", X"77", X"F7", X"7F", X"77", X"7F", X"F7", X"77", X"77", 
X"60", X"88", X"86", X"87", X"88", X"68", X"88", X"86", X"68", X"68", X"67", X"66", X"02", X"80", X"08", X"28", 
X"02", X"06", X"00", X"02", X"60", X"28", X"87", X"88", X"88", X"88", X"88", X"04", X"88", X"80", X"88", X"84", 
X"74", X"7C", X"76", X"67", X"67", X"66", X"74", X"F6", X"67", X"64", X"76", X"67", X"48", X"66", X"48", X"00", 
X"00", X"08", X"00", X"00", X"08", X"08", X"48", X"08", X"08", X"08", X"08", X"08", X"08", X"76", X"54", X"80", 
X"87", X"47", X"48", X"50", X"05", X"00", X"00", X"00", X"80", X"00", X"01", X"00", X"00", X"00", X"00", X"10", 
X"08", X"00", X"00", X"00", X"80", X"01", X"08", X"00", X"00", X"00", X"00", X"50", X"08", X"00", X"08", X"08", 
X"00", X"80", X"00", X"00", X"00", X"00", X"00", X"00", X"01", X"00", X"80", X"00", X"00", X"80", X"00", X"00", 
X"7F", X"6F", X"67", X"7F", X"6F", X"77", X"77", X"78", X"86", X"86", X"88", X"76", X"88", X"86", X"86", X"86", 
X"06", X"86", X"86", X"87", X"68", X"06", X"88", X"86", X"80", X"02", X"08", X"80", X"08", X"08", X"88", X"86", 
X"88", X"47", X"88", X"08", X"84", X"80", X"48", X"68", X"46", X"66", X"47", X"C6", X"6C", X"7C", X"67", X"C7", 
X"C6", X"7C", X"67", X"47", X"66", X"84", X"84", X"00", X"00", X"08", X"08", X"00", X"88", X"80", X"88", X"88", 
X"08", X"80", X"50", X"80", X"40", X"47", X"67", X"40", X"48", X"45", X"67", X"00", X"00", X"00", X"85", X"00", 
X"00", X"80", X"00", X"80", X"08", X"00", X"00", X"08", X"01", X"00", X"80", X"00", X"00", X"80", X"00", X"00", 
X"80", X"08", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"08", X"00", X"80", X"08", X"01", X"08", 
X"00", X"80", X"00", X"80", X"00", X"00", X"50", X"08", X"F7", X"F7", X"76", X"77", X"77", X"76", X"77", X"68", 
X"86", X"88", X"68", X"86", X"76", X"86", X"86", X"88", X"86", X"06", X"86", X"76", X"86", X"02", X"08", X"02", 
X"08", X"00", X"20", X"20", X"02", X"08", X"78", X"80", X"88", X"88", X"80", X"88", X"08", X"08", X"08", X"66", 
X"74", X"74", X"76", X"77", X"67", X"67", X"67", X"66", X"74", X"74", X"76", X"64", X"84", X"86", X"88", X"00", 
X"00", X"08", X"08", X"00", X"80", X"88", X"04", X"88", X"40", X"80", X"80", X"80", X"88", X"44", X"76", X"50", 
X"08", X"74", X"84", X"88", X"08", X"00", X"00", X"80", X"00", X"08", X"00", X"50", X"00", X"00", X"80", X"00", 
X"08", X"00", X"08", X"08", X"00", X"00", X"08", X"00", X"00", X"10", X"00", X"80", X"05", X"08", X"01", X"00", 
X"80", X"10", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"80", X"00", X"00", X"00", 
X"77", X"76", X"77", X"7F", X"6F", X"67", X"76", X"76", X"88", X"67", X"67", X"47", X"67", X"67", X"68", X"66", 
X"76", X"86", X"86", X"86", X"78", X"68", X"00", X"80", X"06", X"08", X"00", X"80", X"20", X"86", X"88", X"60", 
X"88", X"88", X"40", X"80", X"60", X"60", X"64", X"86", X"67", X"46", X"66", X"46", X"7C", X"6C", X"7C", X"7C", 
X"76", X"67", X"47", X"47", X"66", X"68", X"40", X"00", X"00", X"00", X"80", X"80", X"58", X"80", X"88", X"08", 
X"88", X"88", X"04", X"08", X"50", X"87", X"47", X"48", X"45", X"67", X"57", X"04", X"00", X"00", X"00", X"00", 
X"80", X"00", X"00", X"00", X"81", X"00", X"00", X"80", X"00", X"00", X"00", X"00", X"08", X"00", X"00", X"08", 
X"00", X"00", X"80", X"00", X"00", X"00", X"00", X"00", X"00", X"80", X"08", X"01", X"08", X"08", X"08", X"08", 
X"00", X"80", X"80", X"00", X"00", X"80", X"08", X"00", X"7F", X"77", X"77", X"67", X"77", X"67", X"67", X"68", 
X"66", X"74", X"76", X"74", X"74", X"74", X"76", X"76", X"68", X"66", X"86", X"86", X"68", X"86", X"26", X"02", 
X"00", X"06", X"02", X"08", X"00", X"08", X"88", X"06", X"84", X"88", X"80", X"88", X"08", X"08", X"08", X"48", 
X"47", X"47", X"76", X"76", X"67", X"76", X"76", X"67", X"C7", X"66", X"47", X"47", X"48", X"66", X"48", X"80", 
X"00", X"00", X"08", X"00", X"00", X"88", X"88", X"88", X"88", X"08", X"80", X"80", X"08", X"54", X"74", X"80", 
X"04", X"76", X"65", X"88", X"88", X"08", X"00", X"50", X"00", X"00", X"80", X"00", X"00", X"08", X"00", X"00", 
X"80", X"10", X"80", X"00", X"10", X"08", X"00", X"10", X"08", X"00", X"00", X"08", X"00", X"80", X"08", X"08", 
X"00", X"00", X"00", X"80", X"00", X"00", X"00", X"05", X"00", X"00", X"50", X"80", X"10", X"00", X"00", X"00", 
X"76", X"76", X"76", X"F7", X"67", X"67", X"67", X"67", X"67", X"47", X"47", X"47", X"C7", X"47", X"C7", X"47", 
X"47", X"47", X"68", X"68", X"67", X"68", X"00", X"80", X"08", X"00", X"20", X"82", X"00", X"20", X"60", X"80", 
X"88", X"80", X"04", X"06", X"06", X"08", X"48", X"08", X"60", X"84", X"68", X"47", X"6C", X"66", X"67", X"C6", 
X"7C", X"76", X"74", X"66", X"74", X"76", X"80", X"00", X"00", X"00", X"80", X"80", X"88", X"50", X"85", X"78", 
X"48", X"80", X"80", X"50", X"40", X"48", X"47", X"48", X"08", X"47", X"78", X"78", X"80", X"00", X"00", X"00", 
X"80", X"50", X"00", X"08", X"00", X"00", X"00", X"80", X"00", X"00", X"00", X"80", X"00", X"00", X"00", X"00", 
X"00", X"08", X"10", X"00", X"00", X"00", X"00", X"00", X"08", X"01", X"00", X"00", X"81", X"00", X"00", X"00", 
X"00", X"00", X"00", X"00", X"00", X"80", X"08", X"00", X"F7", X"77", X"67", X"77", X"76", X"76", X"76", X"76", 
X"47", X"67", X"C7", X"67", X"47", X"67", X"47", X"47", X"47", X"47", X"66", X"86", X"86", X"76", X"86", X"00", 
X"20", X"00", X"08", X"08", X"00", X"80", X"60", X"60", X"68", X"60", X"08", X"08", X"08", X"80", X"84", X"86", 
X"86", X"80", X"68", X"67", X"67", X"C7", X"66", X"76", X"7C", X"74", X"76", X"76", X"64", X"86", X"48", X"00", 
X"00", X"00", X"08", X"08", X"88", X"77", X"77", X"78", X"88", X"88", X"08", X"08", X"08", X"57", X"47", X"40", 
X"08", X"58", X"40", X"74", X"88", X"80", X"08", X"00", X"00", X"00", X"80", X"00", X"05", X"08", X"01", X"00", 
X"08", X"08", X"00", X"08", X"00", X"50", X"80", X"80", X"80", X"00", X"00", X"80", X"05", X"08", X"00", X"50", 
X"00", X"00", X"80", X"00", X"00", X"05", X"08", X"00", X"80", X"80", X"00", X"08", X"00", X"05", X"00", X"00", 
X"76", X"76", X"77", X"67", X"76", X"76", X"76", X"67", X"47", X"C7", X"67", X"C7", X"6C", X"74", X"7C", X"76", 
X"74", X"74", X"76", X"76", X"68", X"67", X"68", X"00", X"00", X"80", X"20", X"20", X"08", X"08", X"00", X"08", 
X"08", X"00", X"60", X"80", X"40", X"60", X"68", X"68", X"68", X"68", X"40", X"66", X"67", X"66", X"7C", X"76", 
X"67", X"66", X"74", X"67", X"67", X"48", X"60", X"80", X"00", X"00", X"08", X"08", X"88", X"78", X"77", X"85", 
X"08", X"04", X"80", X"80", X"80", X"84", X"75", X"88", X"00", X"08", X"08", X"87", X"88", X"00", X"00", X"08", 
X"00", X"00", X"00", X"80", X"00", X"00", X"00", X"08", X"00", X"00", X"10", X"00", X"00", X"00", X"00", X"00", 
X"05", X"00", X"80", X"10", X"00", X"00", X"00", X"00", X"08", X"00", X"00", X"80", X"00", X"00", X"00", X"00", 
X"00", X"00", X"80", X"00", X"00", X"00", X"08", X"00", X"67", X"77", X"6F", X"67", X"76", X"76", X"76", X"74", 
X"74", X"7C", X"74", X"74", X"77", X"C6", X"74", X"7C", X"74", X"74", X"74", X"76", X"86", X"62", X"86", X"80", 
X"02", X"00", X"00", X"88", X"06", X"88", X"06", X"06", X"06", X"00", X"04", X"08", X"08", X"08", X"06", X"08", 
X"48", X"68", X"84", X"86", X"7C", X"76", X"67", X"47", X"48", X"86", X"74", X"74", X"66", X"68", X"48", X"00", 
X"00", X"00", X"00", X"80", X"88", X"88", X"78", X"88", X"08", X"88", X"08", X"04", X"08", X"84", X"74", X"84", 
X"00", X"00", X"04", X"88", X"48", X"80", X"05", X"00", X"80", X"05", X"00", X"00", X"80", X"00", X"80", X"00", 
X"08", X"00", X"00", X"80", X"08", X"00", X"05", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"08", X"00", 
X"00", X"80", X"00", X"00", X"80", X"80", X"00", X"80", X"05", X"00", X"05", X"08", X"08", X"00", X"00", X"00", 
X"76", X"76", X"77", X"76", X"76", X"76", X"76", X"67", X"47", X"47", X"47", X"C7", X"C6", X"76", X"7C", X"74", 
X"7C", X"74", X"74", X"74", X"76", X"86", X"76", X"80", X"00", X"06", X"00", X"02", X"88", X"80", X"60", X"08", 
X"08", X"06", X"08", X"06", X"04", X"08", X"40", X"86", X"88", X"86", X"86", X"84", X"66", X"7C", X"76", X"67", 
X"68", X"40", X"84", X"08", X"47", X"48", X"60", X"00", X"08", X"00", X"80", X"60", X"80", X"75", X"78", X"88", 
X"80", X"80", X"80", X"80", X"80", X"84", X"74", X"80", X"00", X"50", X"08", X"88", X"78", X"00", X"00", X"00", 
X"00", X"00", X"08", X"00", X"00", X"80", X"00", X"01", X"00", X"08", X"00", X"00", X"00", X"08", X"00", X"00", 
X"08", X"00", X"08", X"08", X"08", X"05", X"00", X"00", X"00", X"00", X"50", X"00", X"00", X"00", X"81", X"00", 
X"00", X"00", X"00", X"00", X"00", X"08", X"08", X"00", X"67", X"76", X"F6", X"77", X"67", X"67", X"67", X"47", 
X"C7", X"67", X"C7", X"47", X"7C", X"74", X"7C", X"76", X"67", X"C7", X"C7", X"64", X"76", X"67", X"67", X"68", 
X"00", X"20", X"80", X"00", X"88", X"80", X"80", X"60", X"60", X"00", X"60", X"00", X"80", X"88", X"00", X"00", 
X"60", X"80", X"86", X"86", X"76", X"67", X"47", X"64", X"84", X"86", X"86", X"86", X"86", X"48", X"66", X"00", 
X"00", X"00", X"00", X"00", X"88", X"78", X"88", X"08", X"48", X"80", X"58", X"08", X"05", X"08", X"88", X"58", 
X"00", X"00", X"04", X"88", X"47", X"08", X"00", X"00", X"80", X"80", X"00", X"08", X"00", X"10", X"08", X"00", 
X"80", X"00", X"08", X"08", X"00", X"00", X"00", X"80", X"00", X"50", X"00", X"00", X"00", X"00", X"00", X"80", 
X"08", X"00", X"00", X"08", X"00", X"00", X"00", X"80", X"00", X"80", X"00", X"00", X"05", X"00", X"00", X"00", 
X"76", X"77", X"67", X"F6", X"76", X"67", X"66", X"74", X"67", X"C7", X"67", X"C7", X"47", X"C7", X"67", X"C7", 
X"47", X"67", X"47", X"67", X"47", X"46", X"76", X"78", X"00", X"00", X"00", X"88", X"86", X"00", X"06", X"00", 
X"00", X"00", X"06", X"04", X"04", X"80", X"04", X"88", X"86", X"80", X"60", X"66", X"47", X"66", X"74", X"68", 
X"68", X"86", X"84", X"86", X"88", X"68", X"48", X"00", X"00", X"00", X"08", X"80", X"08", X"88", X"85", X"88", 
X"08", X"08", X"08", X"04", X"08", X"04", X"08", X"00", X"00", X"00", X"08", X"80", X"84", X"80", X"08", X"00", 
X"00", X"00", X"50", X"01", X"00", X"00", X"00", X"00", X"00", X"80", X"00", X"00", X"08", X"00", X"80", X"00", 
X"00", X"00", X"80", X"01", X"00", X"80", X"00", X"10", X"00", X"08", X"00", X"50", X"08", X"00", X"00", X"00", 
X"80", X"00", X"80", X"08", X"00", X"00", X"50", X"08", X"77", X"67", X"76", X"76", X"76", X"76", X"76", X"67", 
X"47", X"C7", X"47", X"C7", X"67", X"C7", X"C7", X"7C", X"7C", X"76", X"7C", X"74", X"76", X"86", X"67", X"66", 
X"80", X"00", X"20", X"80", X"08", X"60", X"00", X"80", X"48", X"00", X"08", X"00", X"80", X"48", X"00", X"68", 
X"70", X"60", X"88", X"88", X"66", X"76", X"67", X"68", X"68", X"68", X"88", X"86", X"84", X"86", X"86", X"00", 
X"00", X"00", X"00", X"04", X"08", X"88", X"88", X"88", X"88", X"88", X"08", X"08", X"08", X"08", X"08", X"40", 
X"80", X"80", X"00", X"48", X"88", X"80", X"00", X"00", X"50", X"00", X"00", X"00", X"08", X"08", X"08", X"08", 
X"00", X"00", X"05", X"00", X"10", X"00", X"00", X"50", X"08", X"00", X"00", X"08", X"00", X"00", X"80", X"08", 
X"00", X"00", X"00", X"00", X"05", X"00", X"80", X"00", X"00", X"05", X"00", X"00", X"00", X"00", X"00", X"00", 
X"76", X"77", X"6F", X"67", X"76", X"76", X"7C", X"7C", X"66", X"67", X"C7", X"67", X"C7", X"67", X"67", X"C7", 
X"74", X"7C", X"76", X"74", X"74", X"76", X"86", X"76", X"88", X"00", X"08", X"20", X"88", X"00", X"60", X"08", 
X"00", X"00", X"80", X"60", X"68", X"86", X"88", X"06", X"88", X"06", X"84", X"64", X"84", X"67", X"68", X"47", 
X"86", X"87", X"48", X"48", X"68", X"68", X"48", X"00", X"00", X"00", X"00", X"80", X"85", X"88", X"88", X"88", 
X"00", X"80", X"80", X"80", X"80", X"80", X"40", X"80", X"50", X"00", X"08", X"88", X"04", X"80", X"50", X"00", 
X"00", X"80", X"08", X"08", X"00", X"00", X"00", X"01", X"00", X"80", X"00", X"00", X"00", X"80", X"00", X"00", 
X"00", X"05", X"00", X"00", X"08", X"00", X"00", X"00", X"05", X"00", X"80", X"00", X"00", X"00", X"05", X"00", 
X"80", X"00", X"00", X"08", X"00", X"80", X"08", X"00", X"6F", X"67", X"67", X"67", X"67", X"66", X"76", X"7C", 
X"77", X"C6", X"7C", X"76", X"7C", X"7C", X"76", X"7C", X"7C", X"76", X"7C", X"7C", X"74", X"76", X"68", X"68", 
X"62", X"02", X"00", X"00", X"80", X"80", X"06", X"00", X"00", X"00", X"40", X"00", X"04", X"86", X"48", X"68", 
X"68", X"48", X"88", X"68", X"66", X"74", X"76", X"84", X"88", X"88", X"88", X"00", X"68", X"68", X"84", X"80", 
X"00", X"00", X"00", X"00", X"08", X"85", X"80", X"88", X"88", X"04", X"80", X"80", X"50", X"80", X"50", X"80", 
X"00", X"00", X"00", X"88", X"80", X"80", X"00", X"80", X"00", X"00", X"00", X"00", X"00", X"50", X"80", X"00", 
X"01", X"00", X"80", X"08", X"00", X"00", X"80", X"08", X"00", X"00", X"80", X"80", X"00", X"18", X"00", X"80", 
X"00", X"00", X"00", X"80", X"08", X"00", X"00", X"00", X"00", X"00", X"50", X"00", X"00", X"00", X"00", X"00", 
X"77", X"67", X"77", X"66", X"F6", X"76", X"F6", X"67", X"C6", X"7C", X"7C", X"7C", X"77", X"67", X"C7", X"76", 
X"77", X"C7", X"47", X"67", X"66", X"74", X"76", X"76", X"80", X"00", X"02", X"08", X"86", X"00", X"00", X"80", 
X"00", X"00", X"08", X"48", X"68", X"48", X"74", X"86", X"86", X"86", X"84", X"84", X"84", X"66", X"74", X"78", 
X"67", X"78", X"80", X"00", X"48", X"68", X"60", X"00", X"00", X"00", X"00", X"80", X"80", X"88", X"88", X"58", 
X"80", X"80", X"08", X"40", X"80", X"80", X"80", X"80", X"80", X"05", X"00", X"88", X"88", X"08", X"00", X"00", 
X"80", X"08", X"00", X"80", X"00", X"00", X"00", X"80", X"00", X"00", X"00", X"00", X"05", X"00", X"00", X"00", 
X"10", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"80", X"08", X"00", X"00", X"00", X"08", X"00", X"81", 
X"00", X"80", X"00", X"08", X"05", X"08", X"08", X"00", X"76", X"F6", X"6F", X"76", X"67", X"66", X"76", X"76", 
X"7C", X"76", X"7C", X"77", X"C7", X"C7", X"7C", X"7C", X"76", X"7C", X"74", X"7C", X"74", X"76", X"68", X"67", 
X"66", X"02", X"00", X"00", X"08", X"00", X"40", X"06", X"08", X"00", X"00", X"04", X"86", X"74", X"74", X"74", 
X"74", X"74", X"76", X"84", X"76", X"84", X"76", X"67", X"47", X"68", X"08", X"00", X"08", X"48", X"68", X"00", 
X"00", X"00", X"00", X"00", X"88", X"88", X"88", X"87", X"80", X"88", X"00", X"80", X"40", X"80", X"80", X"80", 
X"50", X"00", X"00", X"08", X"40", X"80", X"08", X"00", X"50", X"00", X"50", X"08", X"00", X"08", X"00", X"00", 
X"80", X"08", X"00", X"80", X"00", X"00", X"50", X"08", X"00", X"80", X"00", X"50", X"80", X"05", X"08", X"00", 
X"00", X"05", X"08", X"00", X"50", X"00", X"00", X"00", X"00", X"00", X"80", X"00", X"00", X"00", X"08", X"00", 
X"76", X"77", X"76", X"76", X"F6", X"76", X"F6", X"C7", X"67", X"C7", X"67", X"C7", X"67", X"67", X"C7", X"67", 
X"C7", X"67", X"67", X"67", X"67", X"47", X"66", X"86", X"87", X"80", X"00", X"80", X"80", X"60", X"00", X"00", 
X"00", X"06", X"00", X"06", X"84", X"66", X"76", X"76", X"76", X"76", X"74", X"74", X"84", X"66", X"86", X"78", 
X"74", X"88", X"48", X"48", X"68", X"68", X"84", X"00", X"00", X"00", X"00", X"06", X"08", X"88", X"88", X"77", 
X"50", X"80", X"50", X"80", X"80", X"80", X"85", X"08", X"00", X"00", X"00", X"88", X"88", X"08", X"00", X"00", 
X"00", X"00", X"00", X"00", X"08", X"05", X"00", X"80", X"00", X"01", X"00", X"00", X"80", X"00", X"00", X"00", 
X"00", X"00", X"50", X"00", X"00", X"00", X"00", X"05", X"00", X"00", X"00", X"00", X"00", X"80", X"50", X"08", 
X"00", X"00", X"01", X"00", X"00", X"00", X"00", X"08", X"77", X"66", X"F6", X"74", X"F6", X"67", X"67", X"6F", 
X"66", X"7C", X"F6", X"7C", X"7C", X"76", X"7C", X"76", X"77", X"C7", X"C7", X"C7", X"C7", X"67", X"68", X"68", 
X"66", X"80", X"60", X"08", X"80", X"00", X"08", X"00", X"00", X"00", X"04", X"08", X"47", X"47", X"64", X"74", 
X"74", X"76", X"76", X"84", X"76", X"74", X"74", X"74", X"76", X"84", X"80", X"88", X"84", X"84", X"80", X"00", 
X"00", X"00", X"00", X"00", X"08", X"58", X"88", X"77", X"80", X"80", X"80", X"80", X"80", X"40", X"08", X"08", 
X"08", X"00", X"00", X"00", X"84", X"00", X"08", X"00", X"80", X"08", X"00", X"50", X"00", X"00", X"00", X"00", 
X"08", X"00", X"08", X"00", X"00", X"80", X"80", X"08", X"08", X"00", X"00", X"80", X"08", X"00", X"00", X"00", 
X"08", X"00", X"00", X"80", X"00", X"00", X"00", X"00", X"80", X"80", X"00", X"08", X"08", X"08", X"00", X"00", 
X"76", X"F6", X"76", X"76", X"67", X"6F", X"66", X"C7", X"C7", X"C7", X"6C", X"77", X"C7", X"C7", X"67", X"C7", 
X"C7", X"76", X"77", X"67", X"67", X"47", X"68", X"68", X"68", X"68", X"02", X"06", X"08", X"06", X"00", X"00", 
X"00", X"00", X"00", X"46", X"68", X"46", X"74", X"76", X"76", X"74", X"74", X"86", X"84", X"66", X"67", X"67", 
X"67", X"67", X"64", X"66", X"76", X"86", X"80", X"00", X"00", X"00", X"00", X"00", X"88", X"88", X"88", X"77", 
X"68", X"80", X"80", X"80", X"50", X"80", X"80", X"80", X"80", X"00", X"80", X"08", X"88", X"08", X"00", X"00", 
X"00", X"00", X"00", X"00", X"00", X"08", X"08", X"50", X"00", X"08", X"00", X"10", X"80", X"00", X"00", X"00", 
X"00", X"00", X"00", X"00", X"00", X"08", X"00", X"80", X"00", X"08", X"00", X"00", X"80", X"00", X"80", X"00", 
X"10", X"00", X"80", X"00", X"05", X"00", X"08", X"00", X"76", X"76", X"F7", X"67", X"67", X"66", X"77", X"66", 
X"76", X"7C", X"77", X"C7", X"67", X"7C", X"76", X"77", X"C7", X"C7", X"C7", X"C7", X"68", X"68", X"68", X"68", 
X"62", X"86", X"00", X"80", X"60", X"00", X"08", X"00", X"00", X"60", X"80", X"08", X"64", X"76", X"47", X"66", 
X"47", X"47", X"68", X"47", X"77", X"47", X"64", X"74", X"74", X"76", X"87", X"74", X"74", X"88", X"40", X"00", 
X"00", X"00", X"00", X"08", X"87", X"78", X"87", X"77", X"84", X"80", X"84", X"08", X"08", X"08", X"04", X"08", 
X"05", X"00", X"00", X"00", X"88", X"85", X"08", X"08", X"05", X"08", X"08", X"00", X"80", X"00", X"00", X"00", 
X"80", X"00", X"00", X"00", X"08", X"01", X"08", X"01", X"08", X"08", X"00", X"50", X"80", X"05", X"00", X"00", 
X"05", X"00", X"80", X"01", X"08", X"00", X"08", X"00", X"00", X"00", X"08", X"00", X"00", X"00", X"00", X"80", 
X"76", X"76", X"76", X"76", X"7C", X"7F", X"66", X"F6", X"C7", X"67", X"C7", X"67", X"C7", X"C7", X"7C", X"7C", 
X"77", X"7C", X"77", X"67", X"48", X"86", X"86", X"86", X"86", X"68", X"80", X"88", X"08", X"06", X"00", X"00", 
X"00", X"00", X"40", X"44", X"86", X"47", X"46", X"7C", X"76", X"74", X"74", X"77", X"46", X"74", X"67", X"67", 
X"67", X"47", X"64", X"74", X"76", X"74", X"80", X"00", X"00", X"00", X"00", X"00", X"77", X"77", X"48", X"7F", 
X"88", X"80", X"80", X"80", X"88", X"08", X"08", X"80", X"80", X"00", X"00", X"00", X"07", X"77", X"00", X"00", 
X"00", X"00", X"00", X"10", X"00", X"00", X"00", X"80", X"05", X"00", X"80", X"80", X"00", X"00", X"00", X"08", 
X"00", X"00", X"00", X"00", X"00", X"00", X"08", X"08", X"00", X"00", X"10", X"00", X"00", X"00", X"00", X"08", 
X"08", X"00", X"00", X"08", X"00", X"80", X"50", X"00", X"67", X"6F", X"67", X"66", X"76", X"67", X"C7", X"67", 
X"CF", X"67", X"C7", X"C7", X"C7", X"7C", X"7C", X"77", X"6C", X"77", X"47", X"48", X"48", X"48", X"76", X"78", 
X"68", X"68", X"60", X"80", X"60", X"00", X"00", X"08", X"00", X"00", X"08", X"48", X"68", X"64", X"74", X"67", 
X"C7", X"67", X"68", X"47", X"47", X"67", X"46", X"67", X"C7", X"67", X"47", X"67", X"47", X"48", X"80", X"00", 
X"00", X"00", X"00", X"00", X"77", X"77", X"87", X"77", X"70", X"58", X"08", X"08", X"04", X"80", X"80", X"88", 
X"05", X"08", X"00", X"80", X"06", X"77", X"75", X"08", X"00", X"80", X"08", X"00", X"05", X"08", X"00", X"00", 
X"00", X"00", X"00", X"08", X"00", X"80", X"80", X"00", X"00", X"80", X"80", X"08", X"00", X"80", X"00", X"00", 
X"00", X"00", X"00", X"80", X"50", X"80", X"50", X"00", X"05", X"00", X"80", X"00", X"00", X"00", X"00", X"00", 
X"76", X"76", X"76", X"76", X"76", X"76", X"76", X"C7", X"67", X"C7", X"67", X"67", X"7C", X"77", X"77", X"C7", 
X"C7", X"6C", X"74", X"86", X"86", X"74", X"76", X"86", X"86", X"86", X"88", X"68", X"00", X"60", X"08", X"00", 
X"08", X"00", X"48", X"46", X"48", X"66", X"67", X"47", X"67", X"46", X"84", X"84", X"74", X"74", X"76", X"7C", 
X"76", X"67", X"67", X"47", X"47", X"48", X"00", X"00", X"00", X"00", X"00", X"00", X"77", X"77", X"75", X"7F", 
X"68", X"08", X"05", X"08", X"00", X"80", X"50", X"40", X"80", X"00", X"00", X"00", X"88", X"76", X"7F", X"78", 
X"00", X"05", X"00", X"08", X"00", X"00", X"05", X"00", X"80", X"80", X"00", X"00", X"00", X"00", X"05", X"08", 
X"05", X"00", X"00", X"00", X"50", X"00", X"50", X"00", X"80", X"80", X"88", X"78", X"00", X"00", X"00", X"80", 
X"00", X"00", X"05", X"08", X"08", X"00", X"80", X"80", X"67", X"6F", X"67", X"66", X"6F", X"67", X"67", X"C7", 
X"67", X"6F", X"67", X"66", X"76", X"6C", X"76", X"77", X"C7", X"77", X"67", X"48", X"48", X"74", X"76", X"86", 
X"86", X"76", X"88", X"06", X"80", X"06", X"00", X"00", X"00", X"00", X"04", X"87", X"48", X"47", X"64", X"76", 
X"47", X"47", X"48", X"48", X"66", X"67", X"46", X"76", X"7C", X"7C", X"64", X"74", X"68", X"48", X"48", X"00", 
X"00", X"00", X"00", X"00", X"77", X"77", X"77", X"77", X"78", X"80", X"80", X"80", X"58", X"08", X"08", X"08", 
X"88", X"00", X"50", X"00", X"00", X"77", X"67", X"77", X"78", X"00", X"08", X"00", X"08", X"00", X"00", X"00", 
X"00", X"05", X"80", X"08", X"08", X"00", X"00", X"00", X"00", X"05", X"08", X"00", X"00", X"00", X"08", X"00", 
X"00", X"08", X"77", X"77", X"00", X"80", X"00", X"00", X"00", X"80", X"00", X"00", X"08", X"00", X"00", X"00", 
X"76", X"76", X"76", X"76", X"76", X"67", X"66", X"76", X"C7", X"66", X"67", X"47", X"48", X"76", X"7C", X"76", 
X"7C", X"67", X"47", X"47", X"74", X"88", X"48", X"68", X"68", X"66", X"86", X"88", X"00", X"80", X"00", X"00", 
X"60", X"00", X"68", X"46", X"66", X"48", X"46", X"67", X"C7", X"67", X"46", X"84", X"67", X"46", X"67", X"66", 
X"76", X"76", X"74", X"74", X"74", X"88", X"00", X"00", X"08", X"00", X"00", X"00", X"77", X"77", X"76", X"77", 
X"70", X"84", X"80", X"80", X"80", X"08", X"08", X"80", X"80", X"80", X"00", X"00", X"08", X"47", X"77", X"4F", 
X"77", X"78", X"00", X"00", X"00", X"50", X"08", X"00", X"80", X"00", X"00", X"05", X"00", X"08", X"08", X"00", 
X"08", X"00", X"00", X"08", X"08", X"00", X"00", X"05", X"08", X"77", X"77", X"78", X"00", X"00", X"80", X"80", 
X"80", X"00", X"00", X"80", X"00", X"08", X"08", X"00", X"76", X"F6", X"76", X"67", X"67", X"C7", X"66", X"76", 
X"76", X"74", X"86", X"86", X"84", X"84", X"8C", X"76", X"77", X"C7", X"47", X"47", X"68", X"48", X"00", X"00", 
X"68", X"68", X"68", X"60", X"60", X"08", X"00", X"00", X"00", X"00", X"04", X"88", X"47", X"64", X"74", X"76", 
X"74", X"74", X"76", X"48", X"48", X"67", X"47", X"C7", X"C7", X"47", X"47", X"47", X"68", X"48", X"40", X"00", 
X"00", X"00", X"00", X"00", X"77", X"77", X"77", X"77", X"78", X"80", X"84", X"80", X"84", X"08", X"08", X"05", 
X"08", X"00", X"00", X"50", X"00", X"84", X"77", X"77", X"77", X"77", X"78", X"58", X"00", X"08", X"00", X"05", 
X"08", X"00", X"80", X"00", X"00", X"08", X"00", X"80", X"00", X"00", X"01", X"00", X"00", X"80", X"80", X"87", 
X"77", X"77", X"77", X"58", X"00", X"50", X"00", X"00", X"00", X"08", X"00", X"00", X"08", X"00", X"00", X"80", 
X"76", X"76", X"76", X"76", X"76", X"76", X"67", X"46", X"74", X"77", X"47", X"67", X"48", X"68", X"67", X"47", 
X"C7", X"67", X"47", X"68", X"48", X"00", X"08", X"06", X"06", X"86", X"78", X"88", X"00", X"60", X"00", X"00", 
X"00", X"08", X"48", X"46", X"84", X"86", X"47", X"47", X"47", X"46", X"47", X"67", X"47", X"46", X"67", X"67", 
X"66", X"74", X"67", X"46", X"84", X"88", X"00", X"80", X"00", X"00", X"00", X"00", X"77", X"77", X"77", X"77", 
X"68", X"08", X"80", X"08", X"08", X"08", X"40", X"80", X"88", X"08", X"00", X"00", X"00", X"88", X"7C", X"7C", 
X"77", X"F7", X"F7", X"78", X"08", X"88", X"88", X"88", X"88", X"80", X"80", X"08", X"88", X"88", X"88", X"88", 
X"08", X"08", X"00", X"00", X"50", X"08", X"87", X"77", X"7C", X"77", X"78", X"80", X"00", X"00", X"80", X"50", 
X"08", X"00", X"08", X"08", X"00", X"80", X"80", X"00", X"76", X"F6", X"76", X"66", X"67", X"67", X"66", X"74", 
X"76", X"76", X"74", X"76", X"76", X"74", X"76", X"67", X"C7", X"C7", X"47", X"68", X"86", X"78", X"04", X"08", 
X"86", X"86", X"66", X"66", X"00", X"00", X"08", X"00", X"80", X"00", X"06", X"86", X"66", X"47", X"47", X"64", 
X"74", X"77", X"47", X"47", X"47", X"47", X"6C", X"74", X"74", X"67", X"46", X"74", X"86", X"86", X"00", X"00", 
X"00", X"80", X"00", X"00", X"67", X"77", X"74", X"F7", X"88", X"80", X"88", X"80", X"80", X"80", X"08", X"80", 
X"80", X"50", X"00", X"00", X"00", X"08", X"87", X"74", X"F6", X"57", X"77", X"F7", X"77", X"77", X"77", X"77", 
X"77", X"77", X"77", X"87", X"77", X"77", X"77", X"78", X"80", X"08", X"08", X"00", X"07", X"77", X"7F", X"C7", 
X"77", X"47", X"78", X"08", X"08", X"00", X"00", X"08", X"00", X"08", X"00", X"08", X"00", X"00", X"08", X"00", 
X"76", X"76", X"68", X"77", X"66", X"74", X"67", X"47", X"67", X"C7", X"67", X"47", X"47", X"67", X"47", X"67", 
X"67", X"67", X"47", X"48", X"67", X"68", X"88", X"48", X"68", X"68", X"68", X"88", X"60", X"80", X"00", X"04", 
X"00", X"00", X"68", X"48", X"47", X"46", X"64", X"76", X"74", X"64", X"74", X"66", X"74", X"74", X"76", X"67", 
X"C7", X"66", X"74", X"86", X"84", X"80", X"00", X"00", X"00", X"00", X"00", X"00", X"77", X"77", X"77", X"77", 
X"78", X"50", X"80", X"80", X"80", X"80", X"80", X"48", X"08", X"80", X"00", X"80", X"00", X"08", X"47", X"77", 
X"77", X"F7", X"7F", X"7F", X"7F", X"7F", X"7F", X"7F", X"F7", X"F7", X"F7", X"F7", X"FF", X"FF", X"F7", X"F7", 
X"77", X"77", X"88", X"87", X"77", X"7F", X"77", X"77", X"77", X"77", X"58", X"80", X"00", X"08", X"00", X"00", 
X"08", X"00", X"08", X"00", X"08", X"08", X"00", X"08", X"67", X"67", X"66", X"47", X"67", X"67", X"66", X"7C", 
X"76", X"74", X"76", X"76", X"84", X"76", X"74", X"7C", X"7C", X"74", X"74", X"74", X"88", X"48", X"68", X"86", 
X"86", X"86", X"76", X"68", X"60", X"06", X"00", X"00", X"08", X"00", X"48", X"67", X"48", X"86", X"74", X"74", 
X"74", X"76", X"47", X"47", X"47", X"66", X"47", X"67", X"47", X"47", X"47", X"48", X"68", X"60", X"00", X"00", 
X"00", X"00", X"00", X"00", X"77", X"67", X"77", X"77", X"80", X"84", X"08", X"04", X"05", X"80", X"80", X"80", 
X"80", X"85", X"00", X"00", X"50", X"00", X"87", X"76", X"7C", X"7C", X"77", X"7F", X"7F", X"7F", X"7F", X"7F", 
X"7F", X"7F", X"7F", X"7F", X"77", X"7F", X"7F", X"7F", X"F7", X"F7", X"F7", X"7F", X"CF", X"7C", X"77", X"74", 
X"77", X"77", X"88", X"00", X"50", X"00", X"80", X"80", X"00", X"80", X"00", X"08", X"00", X"50", X"80", X"00", 
X"77", X"67", X"68", X"67", X"47", X"46", X"86", X"76", X"74", X"74", X"74", X"08", X"04", X"84", X"74", X"67", 
X"67", X"C7", X"67", X"47", X"47", X"68", X"47", X"68", X"68", X"68", X"68", X"60", X"80", X"00", X"00", X"80", 
X"00", X"08", X"84", X"68", X"66", X"47", X"46", X"74", X"76", X"84", X"74", X"74", X"64", X"74", X"74", X"66", 
X"74", X"66", X"74", X"68", X"48", X"00", X"00", X"80", X"08", X"00", X"00", X"00", X"77", X"77", X"86", X"77", 
X"48", X"80", X"80", X"80", X"80", X"08", X"08", X"08", X"08", X"80", X"00", X"00", X"00", X"00", X"04", X"87", 
X"77", X"77", X"F7", X"F7", X"F7", X"F7", X"FF", X"7F", X"F7", X"FF", X"7F", X"F7", X"FF", X"7F", X"7F", X"7F", 
X"5F", X"7F", X"7F", X"77", X"77", X"77", X"77", X"77", X"75", X"77", X"80", X"00", X"00", X"00", X"00", X"00", 
X"00", X"00", X"80", X"50", X"00", X"00", X"08", X"00", X"67", X"68", X"68", X"67", X"66", X"76", X"47", X"47", 
X"66", X"84", X"80", X"87", X"08", X"48", X"67", X"47", X"C7", X"47", X"47", X"47", X"47", X"47", X"74", X"76", 
X"86", X"86", X"86", X"86", X"68", X"06", X"00", X"04", X"00", X"00", X"08", X"47", X"47", X"64", X"76", X"48", 
X"44", X"84", X"84", X"84", X"74", X"64", X"74", X"74", X"76", X"84", X"74", X"76", X"86", X"80", X"00", X"00", 
X"00", X"08", X"00", X"00", X"77", X"77", X"77", X"77", X"80", X"80", X"58", X"08", X"08", X"40", X"80", X"50", 
X"80", X"88", X"50", X"00", X"00", X"50", X"08", X"47", X"7C", X"77", X"C7", X"7C", X"F7", X"F7", X"F7", X"F7", 
X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"FF", X"7F", X"7F", X"7F", X"CF", X"7F", X"7C", X"77", X"4F", X"4F", 
X"76", X"78", X"58", X"00", X"80", X"80", X"08", X"08", X"08", X"00", X"00", X"00", X"80", X"80", X"00", X"80", 
X"76", X"66", X"86", X"68", X"67", X"47", X"66", X"74", X"74", X"00", X"84", X"88", X"48", X"86", X"47", X"46", 
X"74", X"7C", X"74", X"74", X"74", X"74", X"47", X"47", X"67", X"68", X"66", X"86", X"00", X"00", X"08", X"00", 
X"08", X"04", X"86", X"68", X"66", X"86", X"67", X"66", X"84", X"84", X"80", X"40", X"84", X"84", X"66", X"74", 
X"64", X"74", X"76", X"84", X"86", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"77", X"77", X"77", X"77", 
X"78", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"80", X"88", X"00", X"00", X"00", X"00", X"88", X"77", 
X"77", X"7F", X"7F", X"7F", X"7F", X"CF", X"7F", X"CF", X"7F", X"7F", X"7F", X"7F", X"7F", X"5F", X"7F", X"7F", 
X"7F", X"77", X"77", X"C7", X"77", X"77", X"77", X"77", X"77", X"70", X"00", X"00", X"00", X"05", X"00", X"00", 
X"00", X"08", X"00", X"80", X"00", X"80", X"80", X"00", X"77", X"86", X"84", X"76", X"66", X"64", X"74", X"74", 
X"88", X"40", X"88", X"48", X"84", X"74", X"76", X"7C", X"74", X"7C", X"74", X"74", X"7C", X"77", X"47", X"47", 
X"66", X"86", X"86", X"86", X"86", X"00", X"40", X"80", X"00", X"00", X"08", X"48", X"47", X"47", X"47", X"47", 
X"48", X"48", X"48", X"40", X"40", X"84", X"84", X"67", X"47", X"66", X"64", X"86", X"86", X"80", X"00", X"00", 
X"00", X"00", X"00", X"00", X"67", X"77", X"77", X"67", X"84", X"80", X"48", X"04", X"08", X"04", X"08", X"04", 
X"80", X"88", X"08", X"08", X"00", X"00", X"00", X"84", X"76", X"76", X"F6", X"F7", X"7F", X"7F", X"7F", X"7F", 
X"CF", X"7F", X"F5", X"F7", X"FF", X"7F", X"7F", X"7F", X"C7", X"F7", X"F7", X"74", X"74", X"7C", X"77", X"77", 
X"77", X"88", X"08", X"00", X"80", X"00", X"00", X"80", X"80", X"08", X"00", X"08", X"00", X"40", X"00", X"80", 
X"66", X"68", X"68", X"67", X"67", X"67", X"46", X"74", X"86", X"88", X"48", X"67", X"47", X"47", X"47", X"47", 
X"47", X"C7", X"47", X"47", X"47", X"C7", X"C7", X"47", X"47", X"68", X"68", X"68", X"60", X"00", X"00", X"60", 
X"00", X"86", X"06", X"68", X"66", X"74", X"67", X"68", X"48", X"84", X"75", X"78", X"50", X"48", X"47", X"47", 
X"66", X"86", X"86", X"86", X"88", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"77", X"77", X"77", X"77", 
X"88", X"08", X"08", X"08", X"08", X"08", X"08", X"80", X"80", X"88", X"80", X"00", X"00", X"00", X"50", X"08", 
X"77", X"7F", X"77", X"F6", X"F6", X"F7", X"F7", X"F7", X"F7", X"F7", X"FF", X"7F", X"C7", X"F7", X"7F", X"77", 
X"F7", X"C7", X"77", X"77", X"77", X"77", X"7C", X"77", X"57", X"08", X"00", X"00", X"08", X"08", X"00", X"00", 
X"00", X"00", X"08", X"00", X"80", X"08", X"00", X"00", X"68", X"68", X"68", X"66", X"47", X"47", X"47", X"47", 
X"68", X"67", X"47", X"47", X"47", X"47", X"C7", X"6C", X"74", X"7C", X"7C", X"74", X"74", X"76", X"7C", X"74", 
X"76", X"86", X"86", X"86", X"86", X"08", X"00", X"00", X"00", X"08", X"08", X"66", X"86", X"67", X"64", X"74", 
X"74", X"76", X"76", X"76", X"77", X"74", X"76", X"74", X"74", X"76", X"86", X"84", X"86", X"00", X"00", X"00", 
X"00", X"00", X"00", X"00", X"77", X"67", X"77", X"77", X"88", X"88", X"80", X"88", X"05", X"08", X"00", X"80", 
X"58", X"88", X"05", X"00", X"80", X"00", X"08", X"08", X"47", X"76", X"F6", X"F7", X"F7", X"F6", X"FC", X"F7", 
X"FF", X"6F", X"6F", X"77", X"F7", X"F7", X"CF", X"7F", X"7F", X"7F", X"C7", X"C7", X"67", X"57", X"77", X"77", 
X"78", X"80", X"00", X"80", X"00", X"08", X"05", X"00", X"80", X"40", X"00", X"80", X"08", X"00", X"80", X"80", 
X"68", X"66", X"86", X"67", X"66", X"74", X"74", X"74", X"74", X"76", X"74", X"74", X"74", X"74", X"7C", X"76", 
X"7C", X"76", X"7C", X"76", X"7C", X"7C", X"77", X"C7", X"47", X"48", X"66", X"86", X"06", X"06", X"06", X"08", 
X"00", X"00", X"84", X"86", X"47", X"48", X"67", X"48", X"47", X"47", X"47", X"C7", X"74", X"77", X"C7", X"74", 
X"74", X"74", X"74", X"80", X"80", X"00", X"00", X"80", X"00", X"80", X"00", X"00", X"77", X"77", X"77", X"76", 
X"88", X"00", X"85", X"08", X"08", X"08", X"50", X"88", X"08", X"08", X"80", X"00", X"00", X"00", X"00", X"08", 
X"77", X"F7", X"F7", X"7C", X"7F", X"6F", X"F7", X"F6", X"F7", X"F7", X"F7", X"F7", X"7F", X"5F", X"77", X"77", 
X"F7", X"77", X"7F", X"77", X"77", X"67", X"77", X"C7", X"78", X"00", X"80", X"00", X"80", X"00", X"00", X"00", 
X"00", X"00", X"80", X"50", X"08", X"08", X"00", X"00", X"66", X"86", X"86", X"84", X"76", X"66", X"47", X"47", 
X"67", X"47", X"67", X"C7", X"C7", X"C7", X"47", X"C7", X"67", X"C7", X"47", X"47", X"47", X"47", X"47", X"47", 
X"47", X"68", X"86", X"86", X"06", X"00", X"00", X"00", X"00", X"06", X"08", X"86", X"74", X"76", X"47", X"67", 
X"4F", X"7C", X"76", X"7C", X"7F", X"C7", X"7C", X"F7", X"67", X"67", X"68", X"60", X"68", X"00", X"00", X"00", 
X"00", X"00", X"00", X"00", X"77", X"76", X"77", X"77", X"84", X"88", X"08", X"08", X"08", X"00", X"80", X"80", 
X"88", X"88", X"88", X"05", X"00", X"80", X"00", X"48", X"67", X"C7", X"6F", X"7F", X"67", X"F6", X"F6", X"FF", 
X"6F", X"CF", X"7C", X"F7", X"F7", X"F7", X"FC", X"F7", X"F6", X"F7", X"77", X"7C", X"7F", X"74", X"77", X"78", 
X"58", X"00", X"50", X"00", X"00", X"80", X"80", X"80", X"08", X"00", X"00", X"08", X"04", X"08", X"08", X"00", 
X"86", X"06", X"86", X"66", X"68", X"47", X"67", X"C7", X"C7", X"C7", X"C7", X"47", X"47", X"C7", X"C7", X"46", 
X"7C", X"74", X"7C", X"74", X"74", X"7C", X"7C", X"7C", X"74", X"74", X"86", X"86", X"88", X"60", X"84", X"00", 
X"00", X"00", X"84", X"84", X"86", X"67", X"67", X"67", X"77", X"C7", X"7C", X"77", X"67", X"7C", X"76", X"7C", 
X"F7", X"47", X"76", X"88", X"80", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"77", X"77", X"77", X"77", 
X"88", X"08", X"08", X"04", X"80", X"84", X"08", X"04", X"80", X"88", X"80", X"00", X"00", X"00", X"08", X"08", 
X"7F", X"7F", X"7F", X"6F", X"7F", X"6F", X"F6", X"F6", X"F7", X"77", X"F7", X"7C", X"7F", X"77", X"F7", X"77", 
X"7F", X"6F", X"6F", X"77", X"76", X"77", X"77", X"77", X"00", X"00", X"00", X"08", X"00", X"00", X"00", X"00", 
X"00", X"00", X"80", X"00", X"08", X"08", X"00", X"80", X"86", X"68", X"68", X"67", X"47", X"47", X"46", X"76", 
X"76", X"76", X"7C", X"7C", X"76", X"7C", X"7C", X"7C", X"74", X"7C", X"7C", X"7C", X"74", X"74", X"74", X"74", 
X"74", X"68", X"68", X"68", X"60", X"60", X"00", X"60", X"80", X"00", X"00", X"86", X"86", X"84", X"76", X"7C", 
X"F6", X"FC", X"7C", X"7C", X"7C", X"76", X"FC", X"77", X"4F", X"77", X"77", X"66", X"76", X"88", X"80", X"88", 
X"68", X"80", X"80", X"00", X"87", X"77", X"87", X"78", X"88", X"84", X"88", X"00", X"80", X"08", X"08", X"80", 
X"80", X"85", X"88", X"00", X"00", X"50", X"00", X"87", X"7F", X"67", X"6F", X"6F", X"6F", X"6F", X"6F", X"F6", 
X"F6", X"F7", X"6F", X"7F", X"77", X"F7", X"7F", X"7F", X"7F", X"77", X"7F", X"6F", X"77", X"77", X"77", X"78", 
X"80", X"80", X"00", X"00", X"80", X"08", X"08", X"05", X"08", X"00", X"00", X"80", X"80", X"80", X"80", X"00", 
X"68", X"68", X"66", X"86", X"66", X"74", X"74", X"7C", X"7C", X"7C", X"76", X"7C", X"7C", X"76", X"7C", X"74", 
X"74", X"74", X"74", X"77", X"47", X"47", X"C7", X"C7", X"47", X"76", X"86", X"86", X"80", X"86", X"00", X"00", 
X"00", X"60", X"86", X"06", X"86", X"77", X"67", X"F7", X"7C", X"77", X"CF", X"67", X"C7", X"6C", X"77", X"FC", 
X"F7", X"C7", X"C7", X"77", X"67", X"76", X"86", X"78", X"87", X"68", X"88", X"00", X"77", X"77", X"76", X"77", 
X"80", X"80", X"08", X"08", X"08", X"80", X"80", X"80", X"85", X"88", X"80", X"80", X"00", X"00", X"05", X"86", 
X"77", X"7F", X"77", X"7F", X"6F", X"7F", X"6F", X"6F", X"F6", X"F6", X"F7", X"77", X"CF", X"77", X"F7", X"CF", 
X"77", X"F6", X"F7", X"77", X"C7", X"7C", X"77", X"78", X"00", X"00", X"80", X"00", X"00", X"00", X"00", X"00", 
X"00", X"08", X"04", X"00", X"80", X"40", X"80", X"08", X"86", X"06", X"86", X"47", X"64", X"7C", X"74", X"74", 
X"76", X"7C", X"7C", X"77", X"C7", X"C7", X"67", X"47", X"47", X"C7", X"C7", X"C7", X"C7", X"47", X"74", X"7C", 
X"74", X"68", X"68", X"68", X"66", X"08", X"08", X"00", X"00", X"00", X"00", X"08", X"47", X"47", X"77", X"CF", 
X"67", X"C7", X"7C", X"F6", X"7C", X"77", X"C7", X"7C", X"7F", X"7F", X"77", X"C7", X"76", X"77", X"77", X"77", 
X"77", X"76", X"86", X"80", X"87", X"78", X"77", X"77", X"48", X"80", X"58", X"05", X"00", X"80", X"50", X"88", 
X"00", X"88", X"58", X"08", X"00", X"00", X"00", X"77", X"C7", X"64", X"76", X"67", X"F6", X"F6", X"F7", X"F6", 
X"F7", X"F6", X"F6", X"F7", X"77", X"F7", X"7F", X"7F", X"C7", X"F7", X"6F", X"77", X"F7", X"77", X"77", X"88", 
X"00", X"00", X"05", X"00", X"80", X"40", X"80", X"08", X"00", X"00", X"00", X"80", X"08", X"80", X"80", X"00", 
X"68", X"68", X"68", X"66", X"74", X"76", X"67", X"C7", X"C7", X"47", X"67", X"C7", X"7C", X"7C", X"7C", X"74", 
X"7C", X"74", X"74", X"76", X"74", X"74", X"47", X"47", X"47", X"76", X"86", X"86", X"08", X"60", X"60", X"80", 
X"00", X"06", X"08", X"86", X"77", X"7F", X"C7", X"7C", X"7C", X"7C", X"76", X"7C", X"76", X"7C", X"76", X"F7", 
X"7C", X"7C", X"7F", X"76", X"FF", X"7C", X"F7", X"CF", X"7F", X"77", X"74", X"80", X"77", X"67", X"78", X"78", 
X"08", X"08", X"00", X"80", X"84", X"08", X"08", X"08", X"08", X"88", X"88", X"00", X"00", X"00", X"08", X"87", 
X"F7", X"F8", X"80", X"86", X"77", X"F6", X"F6", X"F6", X"F6", X"F7", X"76", X"76", X"74", X"77", X"77", X"F7", 
X"F7", X"F7", X"F7", X"F7", X"7F", X"7C", X"F7", X"00", X"08", X"00", X"00", X"00", X"00", X"00", X"00", X"80", 
X"08", X"00", X"00", X"08", X"08", X"08", X"00", X"80", X"86", X"68", X"66", X"86", X"66", X"47", X"47", X"64", 
X"76", X"C7", X"C7", X"C7", X"C7", X"7C", X"74", X"74", X"47", X"47", X"47", X"47", X"47", X"67", X"47", X"47", 
X"44", X"68", X"68", X"68", X"60", X"80", X"00", X"60", X"00", X"00", X"68", X"77", X"7C", X"7F", X"C7", X"C7", 
X"6F", X"67", X"CF", X"67", X"CF", X"67", X"C7", X"6C", X"77", X"FC", X"7C", X"F7", X"C7", X"F7", X"7F", X"C7", 
X"7C", X"74", X"78", X"60", X"87", X"77", X"77", X"77", X"88", X"08", X"40", X"80", X"80", X"80", X"40", X"88", 
X"08", X"08", X"85", X"08", X"00", X"80", X"08", X"76", X"F6", X"76", X"80", X"06", X"F6", X"F7", X"F6", X"F7", 
X"F6", X"76", X"88", X"87", X"04", X"7C", X"F7", X"7F", X"7F", X"77", X"F7", X"7F", X"7F", X"77", X"77", X"80", 
X"50", X"00", X"00", X"00", X"80", X"08", X"00", X"00", X"00", X"00", X"50", X"00", X"80", X"60", X"80", X"00", 
X"68", X"68", X"68", X"47", X"47", X"66", X"67", X"47", X"47", X"47", X"47", X"47", X"C7", X"C7", X"47", X"C7", 
X"44", X"44", X"47", X"44", X"74", X"7C", X"74", X"74", X"77", X"86", X"86", X"86", X"06", X"04", X"08", X"00", 
X"80", X"88", X"77", X"7C", X"F7", X"F6", X"F6", X"F6", X"C7", X"C7", X"66", X"C7", X"67", X"C7", X"67", X"C7", 
X"C7", X"77", X"76", X"F6", X"F7", X"C7", X"C7", X"7F", X"C7", X"7C", X"74", X"00", X"77", X"87", X"87", X"88", 
X"48", X"80", X"80", X"80", X"80", X"80", X"88", X"08", X"88", X"88", X"88", X"80", X"00", X"00", X"86", X"7F", 
X"7F", X"F6", X"F7", X"77", X"77", X"6F", X"6F", X"6F", X"67", X"74", X"08", X"00", X"87", X"7F", X"7C", X"F7", 
X"7F", X"CF", X"7F", X"C7", X"F7", X"F7", X"F7", X"80", X"00", X"80", X"08", X"00", X"00", X"80", X"08", X"08", 
X"08", X"00", X"00", X"80", X"88", X"08", X"00", X"80", X"68", X"68", X"66", X"86", X"47", X"47", X"64", X"7C", 
X"76", X"47", X"C7", X"C7", X"67", X"C7", X"47", X"47", X"74", X"77", X"47", X"47", X"47", X"47", X"47", X"47", 
X"46", X"68", X"60", X"68", X"60", X"60", X"60", X"60", X"08", X"87", X"7F", X"7F", X"C7", X"FC", X"7C", X"F6", 
X"F6", X"7C", X"F7", X"CF", X"67", X"CF", X"6F", X"67", X"6C", X"7C", X"FC", X"77", X"C7", X"77", X"77", X"C7", 
X"7C", X"74", X"78", X"00", X"87", X"78", X"77", X"78", X"80", X"88", X"50", X"80", X"58", X"08", X"05", X"00", 
X"50", X"88", X"88", X"80", X"80", X"00", X"86", X"76", X"F6", X"F6", X"F6", X"76", X"F6", X"F7", X"F6", X"F7", 
X"F6", X"77", X"47", X"47", X"6F", X"6F", X"7F", X"6F", X"77", X"77", X"7F", X"7F", X"77", X"F7", X"77", X"80", 
X"00", X"00", X"00", X"08", X"00", X"00", X"00", X"00", X"08", X"00", X"80", X"00", X"80", X"80", X"80", X"00", 
X"68", X"66", X"86", X"67", X"66", X"74", X"74", X"66", X"7C", X"74", X"67", X"67", X"C7", X"47", X"C7", X"47", 
X"C7", X"C4", X"7C", X"7C", X"74", X"74", X"74", X"74", X"77", X"86", X"86", X"86", X"06", X"00", X"60", X"80", 
X"68", X"7F", X"7F", X"5F", X"77", X"C7", X"6F", X"6C", X"7C", X"76", X"66", X"F6", X"CF", X"67", X"C7", X"C7", 
X"C7", X"6F", X"77", X"C7", X"7C", X"7C", X"74", X"74", X"77", X"47", X"40", X"00", X"78", X"77", X"86", X"78", 
X"84", X"80", X"80", X"40", X"08", X"08", X"08", X"80", X"88", X"88", X"81", X"80", X"00", X"00", X"87", X"77", 
X"6F", X"F6", X"FF", X"F7", X"F6", X"F6", X"F7", X"6F", X"67", X"77", X"77", X"F7", X"F6", X"F7", X"F7", X"F7", 
X"F7", X"F7", X"F7", X"7F", X"7F", X"7F", X"77", X"78", X"00", X"80", X"50", X"00", X"05", X"08", X"05", X"00", 
X"00", X"00", X"08", X"08", X"08", X"40", X"00", X"80", X"68", X"68", X"67", X"64", X"74", X"74", X"74", X"74", 
X"74", X"74", X"74", X"47", X"47", X"47", X"C7", X"47", X"47", X"C7", X"47", X"47", X"47", X"47", X"47", X"47", 
X"44", X"86", X"86", X"86", X"80", X"60", X"00", X"68", X"77", X"CF", X"7F", X"77", X"F6", X"FC", X"76", X"F6", 
X"F6", X"6F", X"7C", X"67", X"66", X"F6", X"76", X"76", X"74", X"7C", X"67", X"C6", X"76", X"74", X"74", X"74", 
X"48", X"68", X"80", X"00", X"76", X"78", X"78", X"78", X"80", X"88", X"80", X"88", X"08", X"04", X"08", X"08", 
X"00", X"88", X"88", X"85", X"08", X"00", X"87", X"6F", X"76", X"F7", X"6F", X"67", X"77", X"6F", X"6F", X"6F", 
X"7F", X"CF", X"6F", X"C7", X"F6", X"F6", X"F7", X"C7", X"77", X"C7", X"7F", X"6F", X"77", X"77", X"F7", X"88", 
X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"08", X"00", X"80", X"00", X"08", X"00", X"80", X"80", X"00", 
X"66", X"86", X"76", X"86", X"66", X"67", X"47", X"47", X"47", X"47", X"C7", X"47", X"C7", X"47", X"47", X"C7", 
X"47", X"47", X"C7", X"47", X"C7", X"44", X"74", X"74", X"76", X"78", X"60", X"60", X"60", X"80", X"60", X"87", 
X"FF", X"7F", X"5F", X"C7", X"C7", X"67", X"CF", X"66", X"7C", X"F4", X"6F", X"6F", X"C7", X"C7", X"CF", X"C6", 
X"7C", X"77", X"76", X"77", X"C7", X"67", X"47", X"47", X"48", X"00", X"00", X"00", X"87", X"78", X"78", X"78", 
X"88", X"40", X"80", X"80", X"80", X"80", X"80", X"80", X"58", X"88", X"88", X"08", X"00", X"00", X"87", X"77", 
X"6F", X"6F", X"6F", X"6F", X"6F", X"76", X"F7", X"7F", X"6F", X"7F", X"6F", X"7F", X"6F", X"77", X"6F", X"7F", 
X"7F", X"7F", X"77", X"7F", X"7F", X"7F", X"57", X"75", X"00", X"00", X"08", X"00", X"80", X"80", X"80", X"00", 
X"00", X"00", X"80", X"00", X"88", X"08", X"00", X"08", X"67", X"66", X"67", X"68", X"67", X"47", X"64", X"76", 
X"47", X"47", X"47", X"64", X"76", X"C7", X"47", X"C7", X"C7", X"47", X"C7", X"47", X"47", X"47", X"44", X"86", 
X"86", X"68", X"68", X"60", X"00", X"60", X"87", X"C7", X"7F", X"7F", X"F7", X"F7", X"77", X"C7", X"67", X"CF", 
X"66", X"F6", X"7C", X"6F", X"6F", X"C7", X"67", X"C7", X"68", X"48", X"68", X"67", X"67", X"46", X"66", X"78", 
X"00", X"06", X"00", X"80", X"88", X"78", X"78", X"76", X"08", X"88", X"80", X"84", X"80", X"80", X"58", X"08", 
X"08", X"88", X"88", X"08", X"08", X"00", X"86", X"F7", X"77", X"F7", X"7F", X"67", X"C7", X"67", X"CF", X"6F", 
X"6F", X"6F", X"6F", X"67", X"F6", X"FF", X"77", X"76", X"77", X"76", X"F7", X"77", X"C7", X"7F", X"77", X"88", 
X"00", X"80", X"00", X"00", X"00", X"00", X"08", X"08", X"08", X"00", X"08", X"00", X"80", X"80", X"80", X"00", 
X"67", X"68", X"66", X"74", X"74", X"74", X"76", X"47", X"C7", X"64", X"7C", X"74", X"67", X"47", X"47", X"47", 
X"47", X"C7", X"47", X"45", X"44", X"54", X"84", X"84", X"76", X"86", X"86", X"80", X"60", X"86", X"87", X"FF", 
X"7D", X"F4", X"F5", X"C7", X"CF", X"66", X"FC", X"76", X"7C", X"6F", X"67", X"6C", X"76", X"F6", X"F4", X"76", 
X"84", X"08", X"48", X"87", X"67", X"67", X"66", X"76", X"08", X"00", X"00", X"00", X"77", X"78", X"87", X"88", 
X"88", X"08", X"05", X"08", X"08", X"08", X"00", X"80", X"85", X"88", X"88", X"80", X"00", X"00", X"87", X"67", 
X"67", X"6F", X"67", X"76", X"77", X"C7", X"67", X"7F", X"6F", X"F7", X"F6", X"FF", X"6F", X"67", X"6F", X"7F", 
X"7F", X"6F", X"7C", X"F7", X"7F", X"77", X"7F", X"88", X"05", X"00", X"08", X"00", X"80", X"40", X"00", X"00", 
X"00", X"00", X"00", X"80", X"60", X"08", X"00", X"80", X"67", X"68", X"67", X"68", X"66", X"47", X"47", X"67", 
X"47", X"47", X"47", X"47", X"47", X"64", X"74", X"7C", X"74", X"74", X"47", X"68", X"77", X"80", X"84", X"84", 
X"76", X"86", X"86", X"60", X"60", X"86", X"77", X"7F", X"7F", X"7F", X"7F", X"7F", X"7C", X"76", X"67", X"C6", 
X"F6", X"7C", X"6F", X"6F", X"7C", X"6C", X"76", X"84", X"86", X"40", X"48", X"67", X"67", X"66", X"76", X"86", 
X"00", X"08", X"06", X"00", X"88", X"77", X"87", X"88", X"88", X"48", X"80", X"80", X"58", X"08", X"40", X"80", 
X"80", X"85", X"88", X"85", X"08", X"00", X"87", X"77", X"77", X"7F", X"6F", X"77", X"47", X"47", X"67", X"6F", 
X"6F", X"6F", X"7F", X"6F", X"6F", X"7F", X"67", X"76", X"77", X"77", X"77", X"77", X"77", X"77", X"77", X"78", 
X"00", X"00", X"00", X"00", X"00", X"08", X"08", X"00", X"80", X"04", X"00", X"00", X"06", X"08", X"00", X"00", 
X"67", X"66", X"86", X"76", X"78", X"67", X"47", X"47", X"47", X"47", X"46", X"74", X"7C", X"74", X"7C", X"74", 
X"45", X"68", X"74", X"78", X"84", X"04", X"04", X"84", X"78", X"68", X"68", X"68", X"68", X"67", X"FF", X"C7", 
X"C7", X"7C", X"F7", X"C7", X"76", X"FC", X"76", X"76", X"F6", X"F6", X"7C", X"7C", X"6F", X"7C", X"76", X"76", 
X"48", X"66", X"84", X"66", X"66", X"F7", X"67", X"68", X"60", X"60", X"00", X"08", X"67", X"86", X"78", X"78", 
X"80", X"00", X"80", X"80", X"80", X"80", X"80", X"88", X"88", X"08", X"88", X"08", X"00", X"08", X"07", X"77", 
X"67", X"67", X"76", X"F6", X"74", X"77", X"7F", X"7F", X"76", X"F6", X"F6", X"77", X"76", X"77", X"77", X"6F", 
X"77", X"F6", X"F7", X"7F", X"6F", X"75", X"F7", X"58", X"00", X"80", X"50", X"00", X"00", X"00", X"00", X"04", 
X"00", X"00", X"08", X"08", X"08", X"00", X"80", X"08", X"67", X"68", X"67", X"67", X"46", X"47", X"47", X"66", 
X"7C", X"74", X"74", X"74", X"74", X"76", X"67", X"47", X"66", X"54", X"80", X"00", X"00", X"04", X"84", X"84", 
X"76", X"86", X"86", X"86", X"67", X"77", X"7F", X"7F", X"7F", X"77", X"F7", X"FF", X"C7", X"6F", X"6C", X"7C", 
X"66", X"CF", X"67", X"6F", X"6F", X"6F", X"C7", X"47", X"47", X"48", X"68", X"67", X"66", X"E6", X"76", X"68", 
X"60", X"00", X"80", X"00", X"87", X"78", X"78", X"84", X"88", X"88", X"08", X"80", X"40", X"80", X"50", X"80", 
X"08", X"88", X"88", X"88", X"08", X"00", X"86", X"77", X"77", X"77", X"77", X"77", X"74", X"7C", X"6F", X"6F", 
X"7F", X"77", X"7F", X"6F", X"77", X"76", X"77", X"77", X"C7", X"76", X"F6", X"77", X"77", X"F7", X"77", X"88", 
X"00", X"00", X"00", X"50", X"80", X"05", X"00", X"00", X"08", X"08", X"00", X"00", X"80", X"80", X"80", X"00", 
X"67", X"66", X"86", X"67", X"88", X"66", X"74", X"74", X"67", X"47", X"C7", X"46", X"74", X"74", X"74", X"84", 
X"84", X"00", X"00", X"04", X"04", X"58", X"48", X"47", X"67", X"68", X"86", X"87", X"7F", X"F7", X"C7", X"7C", 
X"7C", X"7C", X"F7", X"C7", X"C7", X"C7", X"67", X"6F", X"7F", X"67", X"C7", X"C7", X"C7", X"C7", X"6F", X"46", 
X"7C", X"74", X"76", X"67", X"76", X"86", X"67", X"67", X"60", X"80", X"06", X"00", X"88", X"77", X"88", X"88", 
X"08", X"40", X"84", X"08", X"80", X"80", X"80", X"88", X"88", X"85", X"08", X"50", X"80", X"88", X"87", X"76", 
X"76", X"76", X"F6", X"7C", X"77", X"77", X"76", X"F6", X"76", X"F6", X"F7", X"76", X"76", X"F7", X"76", X"F7", 
X"7F", X"77", X"7F", X"7F", X"77", X"77", X"77", X"78", X"10", X"00", X"00", X"00", X"00", X"00", X"08", X"00", 
X"00", X"00", X"08", X"08", X"00", X"80", X"00", X"80", X"76", X"76", X"06", X"86", X"68", X"48", X"64", X"74", 
X"76", X"47", X"64", X"76", X"47", X"47", X"47", X"44", X"80", X"00", X"88", X"08", X"04", X"84", X"84", X"84", 
X"86", X"86", X"86", X"6F", X"7C", X"F7", X"F7", X"77", X"77", X"F5", X"F7", X"F6", X"F6", X"F6", X"F6", X"6C", 
X"66", X"F6", X"F6", X"F6", X"F7", X"FC", X"7C", X"74", X"7C", X"74", X"77", X"66", X"F6", X"76", X"76", X"68", 
X"60", X"60", X"00", X"00", X"88", X"78", X"78", X"88", X"80", X"08", X"08", X"80", X"88", X"08", X"04", X"08", 
X"08", X"88", X"80", X"88", X"05", X"00", X"87", X"77", X"77", X"76", X"77", X"77", X"44", X"76", X"77", X"6F", 
X"77", X"77", X"67", X"77", X"77", X"67", X"77", X"67", X"76", X"7F", X"67", X"6F", X"7F", X"7F", X"97", X"78", 
X"08", X"00", X"00", X"00", X"80", X"80", X"00", X"08", X"00", X"80", X"00", X"08", X"04", X"08", X"00", X"00", 
X"67", X"66", X"86", X"86", X"78", X"68", X"47", X"67", X"47", X"67", X"47", X"47", X"67", X"47", X"66", X"84", 
X"00", X"08", X"48", X"68", X"08", X"84", X"84", X"86", X"76", X"86", X"87", X"7F", X"6F", X"7C", X"7C", X"7C", 
X"7C", X"76", X"FC", X"7C", X"7C", X"66", X"67", X"67", X"6F", X"C6", X"67", X"C6", X"6F", X"6F", X"76", X"7C", 
X"76", X"7C", X"76", X"76", X"67", X"67", X"67", X"76", X"80", X"00", X"80", X"60", X"88", X"87", X"88", X"88", 
X"50", X"88", X"08", X"08", X"04", X"08", X"08", X"08", X"58", X"88", X"88", X"80", X"88", X"08", X"88", X"67", 
X"76", X"77", X"76", X"74", X"77", X"47", X"77", X"76", X"76", X"F6", X"F7", X"67", X"67", X"7F", X"6F", X"7F", 
X"6F", X"77", X"F7", X"F6", X"77", X"F7", X"77", X"78", X"80", X"00", X"80", X"00", X"00", X"00", X"80", X"00", 
X"08", X"00", X"80", X"08", X"00", X"80", X"08", X"00", X"67", X"66", X"06", X"86", X"66", X"84", X"76", X"47", 
X"47", X"C7", X"67", X"47", X"C7", X"47", X"48", X"48", X"48", X"68", X"84", X"78", X"46", X"88", X"84", X"74", 
X"76", X"86", X"67", X"CF", X"5F", X"77", X"7C", X"77", X"77", X"F4", X"7C", X"76", X"F6", X"FC", X"7C", X"F6", 
X"66", X"F6", X"F6", X"FC", X"7C", X"6F", X"C7", X"67", X"C6", X"7C", X"76", X"76", X"76", X"62", X"66", X"86", 
X"76", X"00", X"00", X"00", X"06", X"77", X"88", X"88", X"80", X"80", X"85", X"80", X"80", X"80", X"80", X"80", 
X"08", X"88", X"88", X"50", X"80", X"88", X"07", X"76", X"77", X"76", X"78", X"80", X"58", X"48", X"66", X"77", 
X"77", X"77", X"67", X"77", X"77", X"67", X"76", X"77", X"7F", X"67", X"67", X"F7", X"F7", X"77", X"F7", X"78", 
X"80", X"00", X"00", X"05", X"00", X"50", X"00", X"80", X"00", X"00", X"00", X"08", X"00", X"80", X"08", X"00", 
X"67", X"68", X"60", X"68", X"67", X"68", X"48", X"64", X"74", X"74", X"67", X"46", X"76", X"67", X"47", X"48", 
X"86", X"88", X"68", X"47", X"88", X"48", X"68", X"47", X"47", X"88", X"67", X"77", X"C7", X"CF", X"6F", X"6F", 
X"C7", X"77", X"C7", X"6C", X"7C", X"76", X"67", X"6C", X"F6", X"6F", X"66", X"76", X"F6", X"F6", X"7C", X"76", 
X"77", X"C7", X"67", X"68", X"67", X"66", X"76", X"76", X"00", X"00", X"80", X"08", X"88", X"87", X"88", X"88", 
X"48", X"04", X"80", X"80", X"80", X"80", X"50", X"88", X"88", X"88", X"88", X"88", X"88", X"04", X"88", X"77", 
X"76", X"77", X"84", X"88", X"40", X"50", X"88", X"48", X"67", X"67", X"77", X"67", X"67", X"77", X"77", X"76", 
X"76", X"F7", X"F7", X"67", X"7F", X"7F", X"77", X"78", X"00", X"80", X"00", X"00", X"00", X"00", X"00", X"00", 
X"80", X"08", X"08", X"00", X"80", X"08", X"00", X"00", X"67", X"66", X"60", X"68", X"68", X"67", X"66", X"74", 
X"74", X"67", X"C6", X"74", X"7C", X"74", X"74", X"84", X"74", X"76", X"75", X"74", X"76", X"88", X"84", X"74", 
X"76", X"86", X"7F", X"C7", X"FC", X"76", X"7C", X"77", X"7C", X"77", X"6F", X"67", X"67", X"CF", X"6F", X"67", 
X"67", X"C6", X"FC", X"F6", X"67", X"CF", X"7C", X"76", X"46", X"74", X"86", X"86", X"76", X"86", X"86", X"78", 
X"00", X"00", X"00", X"00", X"88", X"77", X"88", X"88", X"08", X"80", X"84", X"88", X"04", X"08", X"08", X"08", 
X"08", X"88", X"80", X"80", X"50", X"80", X"87", X"67", X"77", X"67", X"78", X"88", X"88", X"47", X"48", X"88", 
X"88", X"87", X"67", X"87", X"67", X"67", X"67", X"6F", X"77", X"76", X"77", X"F7", X"77", X"77", X"77", X"78", 
X"05", X"00", X"80", X"00", X"00", X"80", X"50", X"80", X"00", X"00", X"00", X"80", X"08", X"00", X"80", X"80", 
X"67", X"68", X"66", X"60", X"66", X"86", X"74", X"66", X"74", X"74", X"76", X"74", X"76", X"76", X"74", X"78", 
X"77", X"47", X"68", X"67", X"57", X"67", X"48", X"47", X"47", X"67", X"7C", X"76", X"F7", X"6F", X"67", X"7C", 
X"77", X"7C", X"74", X"7C", X"76", X"66", X"C7", X"6F", X"6F", X"6F", X"67", X"67", X"C7", X"67", X"C7", X"C7", 
X"74", X"74", X"76", X"00", X"06", X"26", X"F6", X"76", X"08", X"00", X"06", X"00", X"88", X"87", X"88", X"88", 
X"88", X"88", X"08", X"08", X"08", X"08", X"04", X"08", X"88", X"58", X"88", X"88", X"88", X"08", X"87", X"77", 
X"67", X"77", X"67", X"48", X"67", X"78", X"56", X"74", X"86", X"88", X"88", X"67", X"77", X"77", X"7F", X"67", 
X"6F", X"7F", X"6F", X"6F", X"77", X"7F", X"57", X"78", X"80", X"00", X"00", X"80", X"00", X"00", X"00", X"05", 
X"08", X"00", X"40", X"08", X"00", X"80", X"00", X"00", X"66", X"68", X"68", X"68", X"68", X"66", X"76", X"86", 
X"47", X"47", X"C7", X"66", X"C7", X"64", X"74", X"64", X"47", X"87", X"47", X"47", X"67", X"67", X"74", X"74", 
X"86", X"8C", X"7F", X"7C", X"7C", X"7C", X"76", X"F6", X"FC", X"77", X"67", X"66", X"F6", X"F7", X"C7", X"66", 
X"C7", X"66", X"FC", X"F6", X"7C", X"F6", X"F6", X"74", X"76", X"86", X"08", X"00", X"00", X"87", X"67", X"08", 
X"00", X"00", X"00", X"00", X"88", X"77", X"70", X"88", X"08", X"08", X"80", X"80", X"80", X"80", X"88", X"08", 
X"80", X"88", X"80", X"80", X"88", X"00", X"86", X"77", X"F6", X"77", X"77", X"77", X"76", X"76", X"74", X"78", 
X"77", X"76", X"78", X"77", X"67", X"67", X"67", X"F7", X"76", X"77", X"77", X"77", X"77", X"7F", X"79", X"78", 
X"00", X"00", X"00", X"00", X"80", X"08", X"00", X"00", X"00", X"00", X"00", X"04", X"00", X"80", X"08", X"00", 
X"76", X"76", X"68", X"66", X"06", X"86", X"86", X"67", X"46", X"66", X"67", X"47", X"67", X"C7", X"67", X"88", 
X"74", X"74", X"77", X"47", X"C7", X"77", X"67", X"44", X"74", X"77", X"C7", X"C7", X"77", X"76", X"76", X"77", 
X"67", X"7C", X"F6", X"7C", X"67", X"66", X"F6", X"F6", X"76", X"F6", X"67", X"6F", X"66", X"7C", X"7C", X"7C", 
X"74", X"88", X"00", X"00", X"00", X"00", X"86", X"00", X"08", X"00", X"00", X"00", X"88", X"77", X"75", X"88", 
X"40", X"88", X"08", X"40", X"80", X"80", X"80", X"88", X"88", X"88", X"58", X"88", X"50", X"80", X"87", X"76", 
X"77", X"76", X"77", X"67", X"67", X"77", X"77", X"47", X"47", X"77", X"67", X"67", X"77", X"F6", X"F6", X"76", 
X"F7", X"6F", X"6F", X"6F", X"77", X"77", X"77", X"78", X"08", X"05", X"00", X"50", X"00", X"00", X"08", X"00", 
X"80", X"80", X"80", X"00", X"80", X"00", X"80", X"00", X"68", X"68", X"66", X"86", X"68", X"66", X"67", X"68", 
X"67", X"47", X"47", X"47", X"47", X"67", X"44", X"47", X"65", X"7C", X"76", X"57", X"47", X"47", X"76", X"54", 
X"74", X"F7", X"F6", X"F6", X"C7", X"C7", X"7C", X"76", X"F6", X"76", X"76", X"76", X"7C", X"76", X"6C", X"7C", 
X"F6", X"6F", X"C7", X"C7", X"C7", X"67", X"C7", X"67", X"68", X"40", X"08", X"00", X"80", X"00", X"00", X"06", 
X"00", X"00", X"00", X"00", X"88", X"77", X"78", X"80", X"88", X"08", X"80", X"88", X"05", X"80", X"84", X"08", 
X"08", X"88", X"80", X"80", X"88", X"80", X"88", X"77", X"67", X"77", X"78", X"77", X"67", X"67", X"67", X"77", 
X"76", X"77", X"77", X"76", X"76", X"77", X"7F", X"6F", X"67", X"77", X"77", X"77", X"77", X"77", X"77", X"88", 
X"00", X"00", X"00", X"00", X"00", X"50", X"00", X"00", X"00", X"00", X"80", X"80", X"08", X"00", X"00", X"80", 
X"67", X"66", X"86", X"86", X"66", X"86", X"84", X"67", X"48", X"46", X"74", X"67", X"47", X"C7", X"67", X"47", 
X"76", X"74", X"7C", X"7C", X"74", X"76", X"F4", X"74", X"76", X"7C", X"7C", X"76", X"F6", X"76", X"F6", X"76", 
X"76", X"76", X"76", X"67", X"67", X"C7", X"F6", X"76", X"6F", X"67", X"6F", X"67", X"67", X"C7", X"7C", X"76", 
X"78", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"08", X"00", X"00", X"00", X"88", X"87", X"78", X"88", 
X"05", X"08", X"88", X"04", X"00", X"80", X"80", X"88", X"88", X"88", X"88", X"88", X"80", X"80", X"88", X"67", 
X"77", X"67", X"67", X"77", X"77", X"76", X"76", X"76", X"77", X"86", X"87", X"87", X"77", X"6F", X"67", X"77", 
X"7F", X"67", X"67", X"77", X"77", X"77", X"79", X"80", X"00", X"00", X"00", X"80", X"00", X"00", X"80", X"80", 
X"00", X"00", X"00", X"08", X"00", X"80", X"80", X"00", X"62", X"68", X"68", X"68", X"86", X"66", X"68", X"66", 
X"76", X"74", X"67", X"47", X"66", X"74", X"74", X"76", X"47", X"74", X"74", X"74", X"47", X"47", X"74", X"47", 
X"C7", X"F6", X"F7", X"C7", X"67", X"66", X"76", X"7C", X"76", X"7C", X"76", X"76", X"67", X"66", X"67", X"C7", 
X"67", X"CF", X"66", X"FC", X"76", X"76", X"67", X"48", X"60", X"08", X"08", X"08", X"08", X"08", X"00", X"80", 
X"00", X"08", X"00", X"00", X"08", X"77", X"75", X"80", X"80", X"48", X"08", X"08", X"80", X"80", X"80", X"50", 
X"88", X"08", X"88", X"80", X"50", X"40", X"08", X"77", X"77", X"77", X"76", X"86", X"74", X"77", X"77", X"76", 
X"78", X"78", X"67", X"67", X"67", X"77", X"6F", X"67", X"67", X"7F", X"7C", X"77", X"77", X"77", X"77", X"85", 
X"80", X"80", X"00", X"08", X"08", X"00", X"00", X"50", X"08", X"00", X"08", X"00", X"05", X"00", X"00", X"00", 
X"86", X"86", X"86", X"06", X"68", X"86", X"86", X"86", X"68", X"67", X"46", X"74", X"74", X"76", X"47", X"47", 
X"47", X"77", X"74", X"77", X"74", X"F7", X"67", X"47", X"7C", X"7C", X"76", X"76", X"F6", X"76", X"76", X"76", 
X"76", X"76", X"84", X"86", X"66", X"7C", X"F6", X"7C", X"76", X"66", X"7C", X"76", X"74", X"74", X"76", X"78", 
X"00", X"80", X"00", X"00", X"00", X"00", X"08", X"00", X"08", X"00", X"00", X"00", X"05", X"87", X"78", X"88", 
X"80", X"80", X"80", X"80", X"08", X"40", X"88", X"88", X"85", X"88", X"50", X"88", X"80", X"88", X"50", X"86", 
X"76", X"77", X"67", X"77", X"87", X"84", X"88", X"88", X"84", X"88", X"87", X"76", X"F6", X"F6", X"77", X"7F", 
X"6F", X"67", X"77", X"77", X"77", X"77", X"77", X"78", X"80", X"00", X"00", X"00", X"00", X"05", X"00", X"00", 
X"00", X"08", X"00", X"50", X"00", X"08", X"08", X"00", X"68", X"68", X"68", X"67", X"67", X"68", X"66", X"68", 
X"66", X"84", X"76", X"66", X"47", X"C7", X"47", X"47", X"C7", X"C7", X"76", X"7C", X"76", X"76", X"54", X"7C", 
X"7F", X"67", X"CF", X"64", X"7C", X"7C", X"76", X"76", X"74", X"86", X"84", X"88", X"66", X"76", X"66", X"6F", 
X"6F", X"C7", X"67", X"C7", X"64", X"76", X"84", X"86", X"00", X"00", X"00", X"00", X"60", X"80", X"00", X"80", 
X"00", X"00", X"00", X"00", X"08", X"87", X"78", X"80", X"88", X"08", X"80", X"88", X"00", X"80", X"00", X"80", 
X"80", X"80", X"88", X"08", X"08", X"00", X"08", X"88", X"77", X"87", X"88", X"88", X"88", X"88", X"88", X"48", 
X"88", X"88", X"08", X"88", X"88", X"88", X"68", X"68", X"88", X"88", X"78", X"77", X"75", X"88", X"88", X"88", 
X"85", X"08", X"05", X"08", X"00", X"00", X"00", X"80", X"05", X"00", X"00", X"00", X"80", X"05", X"00", X"00", 
X"76", X"86", X"86", X"76", X"67", X"66", X"86", X"86", X"86", X"68", X"68", X"47", X"68", X"67", X"44", X"74", 
X"74", X"76", X"77", X"77", X"47", X"47", X"67", X"7F", X"C7", X"FC", X"76", X"7C", X"76", X"76", X"74", X"74", 
X"86", X"86", X"88", X"04", X"86", X"67", X"6F", X"66", X"76", X"76", X"67", X"66", X"86", X"84", X"88", X"00", 
X"08", X"08", X"06", X"00", X"00", X"00", X"00", X"00", X"06", X"00", X"80", X"00", X"08", X"87", X"88", X"80", 
X"80", X"40", X"50", X"05", X"08", X"05", X"00", X"00", X"00", X"00", X"00", X"00", X"05", X"08", X"08", X"48", 
X"08", X"06", X"08", X"04", X"00", X"84", X"08", X"08", X"00", X"08", X"08", X"08", X"06", X"88", X"88", X"08", 
X"88", X"68", X"86", X"88", X"88", X"88", X"88", X"80", X"00", X"00", X"00", X"00", X"00", X"80", X"00", X"00", 
X"00", X"00", X"80", X"80", X"00", X"00", X"08", X"00", X"76", X"77", X"26", X"77", X"E7", X"66", X"86", X"66", 
X"86", X"86", X"48", X"47", X"64", X"76", X"74", X"74", X"47", X"C7", X"C4", X"C7", X"65", X"C7", X"C7", X"6F", 
X"C7", X"67", X"C6", X"76", X"74", X"76", X"74", X"76", X"68", X"60", X"40", X"00", X"04", X"76", X"67", X"C7", 
X"C7", X"C7", X"66", X"84", X"84", X"86", X"06", X"00", X"00", X"00", X"00", X"00", X"00", X"08", X"00", X"80", 
X"00", X"00", X"00", X"00", X"08", X"87", X"88", X"50", X"80", X"00", X"00", X"00", X"00", X"00", X"08", X"08", 
X"08", X"00", X"50", X"00", X"00", X"00", X"88", X"88", X"68", X"78", X"77", X"77", X"77", X"77", X"77", X"87", 
X"86", X"88", X"68", X"68", X"80", X"80", X"88", X"86", X"88", X"88", X"88", X"88", X"88", X"88", X"88", X"80", 
X"80", X"08", X"00", X"05", X"00", X"08", X"05", X"08", X"08", X"00", X"00", X"05", X"08", X"00", X"08", X"00", 
X"76", X"76", X"7F", X"66", X"76", X"67", X"66", X"86", X"66", X"86", X"86", X"68", X"47", X"47", X"C7", X"47", 
X"44", X"84", X"77", X"45", X"67", X"47", X"7F", X"C7", X"7C", X"F6", X"77", X"C7", X"67", X"C7", X"47", X"67", 
X"48", X"80", X"60", X"00", X"08", X"48", X"67", X"67", X"67", X"67", X"47", X"48", X"48", X"60", X"00", X"00", 
X"80", X"08", X"00", X"80", X"80", X"06", X"00", X"00", X"80", X"00", X"00", X"00", X"08", X"18", X"88", X"00", 
X"00", X"80", X"80", X"80", X"08", X"08", X"00", X"05", X"00", X"00", X"00", X"00", X"08", X"87", X"7F", X"7F", 
X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"FF", X"7F", X"7F", X"7F", X"7F", X"7F", X"6F", X"77", 
X"F7", X"7F", X"77", X"7F", X"7F", X"77", X"78", X"88", X"88", X"00", X"80", X"00", X"00", X"00", X"00", X"00", 
X"00", X"50", X"00", X"00", X"00", X"08", X"00", X"08", X"67", X"6F", X"66", X"7E", X"67", X"66", X"86", X"86", 
X"86", X"86", X"68", X"48", X"66", X"67", X"67", X"47", X"47", X"45", X"44", X"74", X"74", X"7C", X"77", X"FC", 
X"76", X"7C", X"76", X"7C", X"76", X"7C", X"74", X"86", X"84", X"60", X"00", X"80", X"00", X"84", X"76", X"67", 
X"C7", X"67", X"48", X"68", X"60", X"80", X"00", X"00", X"00", X"08", X"00", X"00", X"00", X"00", X"00", X"00", 
X"00", X"80", X"80", X"00", X"08", X"88", X"88", X"80", X"50", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
X"08", X"00", X"80", X"07", X"77", X"FF", X"7F", X"7F", X"7F", X"F7", X"F7", X"F7", X"FF", X"7F", X"7F", X"CF", 
X"7F", X"7F", X"7F", X"7E", X"F6", X"FF", X"7F", X"F7", X"F6", X"F7", X"FF", X"F7", X"F7", X"FF", X"F7", X"FF", 
X"7F", X"7F", X"77", X"F7", X"77", X"78", X"88", X"80", X"00", X"05", X"08", X"08", X"00", X"10", X"00", X"00", 
X"76", X"E6", X"7F", X"67", X"67", X"62", X"66", X"86", X"66", X"68", X"68", X"68", X"48", X"64", X"76", X"76", 
X"84", X"76", X"84", X"47", X"47", X"F7", X"FC", X"77", X"CF", X"6F", X"66", X"76", X"7C", X"76", X"74", X"68", 
X"60", X"08", X"40", X"06", X"04", X"06", X"84", X"76", X"76", X"74", X"86", X"84", X"86", X"00", X"08", X"00", 
X"60", X"00", X"00", X"08", X"00", X"08", X"00", X"80", X"00", X"00", X"00", X"00", X"80", X"80", X"80", X"80", 
X"00", X"85", X"00", X"50", X"80", X"50", X"08", X"00", X"00", X"00", X"05", X"7F", X"7F", X"7F", X"F7", X"F7", 
X"F7", X"FF", X"7F", X"F6", X"F7", X"FC", X"F7", X"F7", X"F7", X"F6", X"FF", X"7F", X"7F", X"F6", X"F6", X"FF", 
X"FF", X"7F", X"6F", X"6F", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"FF", X"7F", X"FF", X"7F", X"F7", X"F7", 
X"F7", X"88", X"00", X"01", X"00", X"08", X"08", X"00", X"76", X"76", X"66", X"6E", X"76", X"68", X"68", X"60", 
X"86", X"76", X"66", X"86", X"84", X"86", X"47", X"67", X"47", X"47", X"47", X"74", X"7C", X"76", X"F6", X"F6", 
X"76", X"6F", X"C7", X"C6", X"76", X"76", X"76", X"86", X"86", X"00", X"00", X"00", X"00", X"04", X"86", X"48", 
X"64", X"86", X"84", X"86", X"08", X"00", X"00", X"00", X"00", X"00", X"80", X"00", X"80", X"00", X"00", X"00", 
X"00", X"00", X"00", X"00", X"00", X"88", X"50", X"80", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"80", 
X"05", X"08", X"77", X"F7", X"FF", X"5F", X"7F", X"FF", X"7F", X"7F", X"6F", X"F7", X"FF", X"7F", X"F7", X"FF", 
X"6F", X"FF", X"6F", X"6F", X"F6", X"FF", X"F7", X"F6", X"7F", X"6F", X"FF", X"7F", X"7F", X"7F", X"7F", X"7F", 
X"7F", X"F7", X"F7", X"F7", X"7F", X"F7", X"FF", X"7F", X"7F", X"7F", X"77", X"88", X"08", X"00", X"00", X"00", 
X"67", X"67", X"F6", X"77", X"67", X"66", X"86", X"60", X"68", X"68", X"68", X"68", X"60", X"48", X"64", X"76", 
X"74", X"74", X"74", X"77", X"F7", X"FC", X"77", X"C7", X"CF", X"67", X"67", X"7C", X"7C", X"76", X"74", X"88", 
X"00", X"06", X"06", X"00", X"84", X"06", X"84", X"84", X"86", X"84", X"86", X"86", X"86", X"00", X"08", X"00", 
X"80", X"00", X"06", X"00", X"00", X"06", X"00", X"06", X"00", X"00", X"00", X"00", X"80", X"80", X"88", X"05", 
X"00", X"08", X"08", X"00", X"80", X"08", X"05", X"00", X"00", X"87", X"F9", X"F7", X"F7", X"77", X"7F", X"7F", 
X"7F", X"7F", X"F7", X"FF", X"6F", X"F7", X"F7", X"F7", X"FF", X"7F", X"FF", X"F7", X"FF", X"7E", X"7F", X"FF", 
X"FF", X"F7", X"6F", X"F6", X"F6", X"FF", X"6F", X"F6", X"F6", X"FF", X"6F", X"F6", X"F7", X"F7", X"7F", X"7F", 
X"F7", X"F7", X"FF", X"77", X"80", X"80", X"50", X"80", X"67", X"66", X"76", X"76", X"76", X"76", X"06", X"86", 
X"86", X"86", X"66", X"68", X"68", X"48", X"47", X"47", X"C7", X"67", X"C7", X"C7", X"C7", X"7F", X"6F", X"C7", 
X"4F", X"6F", X"C6", X"F6", X"77", X"47", X"68", X"40", X"68", X"00", X"00", X"00", X"06", X"00", X"86", X"84", 
X"06", X"68", X"48", X"60", X"00", X"00", X"00", X"00", X"00", X"80", X"00", X"00", X"80", X"00", X"00", X"00", 
X"00", X"08", X"00", X"00", X"50", X"80", X"08", X"00", X"08", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
X"88", X"9F", X"7F", X"9F", X"78", X"00", X"08", X"88", X"04", X"07", X"77", X"FF", X"7F", X"7F", X"7F", X"F7", 
X"F6", X"F7", X"F6", X"F7", X"E7", X"F7", X"F6", X"F6", X"F6", X"FF", X"F6", X"FF", X"FF", X"6F", X"F7", X"FF", 
X"F7", X"FF", X"6F", X"FF", X"77", X"67", X"67", X"7F", X"7F", X"7F", X"7F", X"7F", X"F8", X"00", X"00", X"00", 
X"76", X"76", X"76", X"76", X"76", X"86", X"86", X"06", X"06", X"76", X"76", X"86", X"86", X"86", X"04", X"86", 
X"76", X"74", X"77", X"6F", X"7C", X"F4", X"F6", X"76", X"FC", X"76", X"77", X"C7", X"C7", X"68", X"48", X"80", 
X"00", X"60", X"60", X"60", X"00", X"44", X"04", X"86", X"04", X"86", X"86", X"04", X"80", X"00", X"08", X"00", 
X"80", X"00", X"08", X"06", X"00", X"08", X"00", X"00", X"08", X"00", X"00", X"00", X"08", X"08", X"08", X"08", 
X"00", X"50", X"08", X"50", X"05", X"00", X"08", X"00", X"77", X"77", X"7F", X"77", X"78", X"00", X"00", X"00", 
X"00", X"80", X"47", X"F7", X"FF", X"6F", X"F7", X"FF", X"7F", X"F6", X"FF", X"7F", X"7F", X"F6", X"FF", X"7F", 
X"FF", X"6F", X"7F", X"7F", X"6F", X"F7", X"6F", X"6F", X"7F", X"6F", X"F7", X"F6", X"62", X"82", X"7F", X"F6", 
X"F7", X"F7", X"F7", X"F7", X"7F", X"80", X"80", X"80", X"86", X"88", X"67", X"67", X"68", X"26", X"86", X"82", 
X"68", X"67", X"67", X"66", X"84", X"06", X"84", X"84", X"74", X"74", X"7C", X"7F", X"77", X"7C", X"6F", X"C7", 
X"67", X"CF", X"6F", X"67", X"67", X"68", X"86", X"06", X"00", X"00", X"00", X"00", X"40", X"00", X"60", X"48", 
X"40", X"64", X"86", X"80", X"60", X"00", X"00", X"00", X"60", X"80", X"00", X"00", X"80", X"00", X"08", X"00", 
X"00", X"00", X"00", X"00", X"00", X"50", X"80", X"50", X"00", X"00", X"00", X"00", X"00", X"80", X"00", X"07", 
X"7F", X"9F", X"97", X"F9", X"88", X"08", X"00", X"88", X"00", X"00", X"00", X"67", X"7F", X"F7", X"FF", X"6F", 
X"F7", X"FF", X"7F", X"F6", X"F7", X"FF", X"6F", X"7E", X"7F", X"F7", X"FE", X"7F", X"F6", X"FF", X"FF", X"F6", 
X"F7", X"72", X"67", X"77", X"36", X"77", X"67", X"F7", X"F7", X"F7", X"F7", X"7F", X"7F", X"90", X"80", X"00", 
X"88", X"68", X"86", X"82", X"68", X"68", X"68", X"68", X"68", X"67", X"66", X"76", X"86", X"06", X"06", X"04", 
X"84", X"76", X"7F", X"7C", X"7C", X"F7", X"67", X"6F", X"CF", X"67", X"C7", X"C7", X"67", X"48", X"60", X"00", 
X"80", X"60", X"84", X"08", X"06", X"04", X"86", X"06", X"04", X"86", X"06", X"00", X"80", X"08", X"00", X"00", 
X"00", X"00", X"08", X"00", X"08", X"08", X"00", X"00", X"00", X"00", X"80", X"00", X"80", X"00", X"88", X"00", 
X"80", X"80", X"00", X"80", X"00", X"08", X"08", X"79", X"77", X"F7", X"7F", X"7F", X"80", X"00", X"50", X"00", 
X"00", X"08", X"00", X"80", X"77", X"77", X"6F", X"77", X"7F", X"6F", X"7F", X"7F", X"F6", X"FF", X"F7", X"F7", 
X"F6", X"FE", X"7F", X"7F", X"7F", X"F6", X"F6", X"72", X"62", X"86", X"22", X"62", X"28", X"28", X"28", X"7F", 
X"6F", X"7F", X"7F", X"77", X"F7", X"78", X"00", X"88", X"88", X"68", X"06", X"88", X"68", X"60", X"68", X"68", 
X"26", X"76", X"76", X"86", X"86", X"04", X"86", X"06", X"84", X"77", X"C7", X"7F", X"7C", X"7C", X"FC", X"76", 
X"76", X"F6", X"7F", X"C7", X"76", X"88", X"08", X"04", X"00", X"00", X"00", X"40", X"08", X"00", X"48", X"40", 
X"68", X"48", X"48", X"60", X"60", X"00", X"00", X"80", X"00", X"80", X"06", X"80", X"06", X"00", X"08", X"00", 
X"80", X"00", X"00", X"00", X"08", X"80", X"08", X"00", X"00", X"08", X"00", X"00", X"80", X"00", X"07", X"7F", 
X"79", X"7F", X"97", X"9F", X"58", X"00", X"00", X"00", X"85", X"00", X"00", X"80", X"86", X"77", X"77", X"E7", 
X"6F", X"67", X"E7", X"77", X"F7", X"F6", X"FF", X"6F", X"FF", X"7F", X"7F", X"7F", X"E7", X"F7", X"28", X"28", 
X"88", X"28", X"72", X"87", X"67", X"28", X"6F", X"7F", X"F7", X"F6", X"F7", X"F7", X"7F", X"78", X"10", X"87", 
X"08", X"88", X"60", X"86", X"86", X"86", X"88", X"68", X"67", X"67", X"67", X"67", X"68", X"60", X"48", X"68", 
X"68", X"67", X"F7", X"C7", X"77", X"6F", X"67", X"CF", X"C7", X"CF", X"67", X"76", X"74", X"86", X"00", X"00", 
X"80", X"80", X"00", X"00", X"40", X"40", X"60", X"60", X"40", X"68", X"68", X"08", X"80", X"06", X"00", X"00", 
X"60", X"00", X"00", X"00", X"80", X"08", X"00", X"00", X"00", X"00", X"00", X"00", X"80", X"08", X"88", X"05", 
X"00", X"50", X"08", X"00", X"00", X"80", X"87", X"97", X"F7", X"79", X"F7", X"77", X"F0", X"80", X"80", X"00", 
X"00", X"08", X"50", X"00", X"88", X"77", X"67", X"76", X"72", X"77", X"77", X"6F", X"FF", X"FF", X"7F", X"F7", 
X"F6", X"FF", X"6F", X"F7", X"77", X"26", X"72", X"72", X"62", X"82", X"76", X"27", X"27", X"63", X"27", X"F7", 
X"F6", X"F7", X"F7", X"7F", X"7F", X"77", X"00", X"7F", X"60", X"80", X"60", X"08", X"86", X"28", X"66", X"86", 
X"86", X"27", X"67", X"68", X"68", X"48", X"40", X"48", X"67", X"77", X"C7", X"7F", X"C7", X"C7", X"C7", X"6F", 
X"67", X"7C", X"7C", X"76", X"78", X"80", X"00", X"40", X"00", X"40", X"60", X"80", X"00", X"40", X"04", X"84", 
X"86", X"04", X"84", X"06", X"80", X"00", X"80", X"00", X"80", X"80", X"06", X"00", X"80", X"00", X"60", X"80", 
X"06", X"08", X"08", X"00", X"85", X"88", X"88", X"00", X"00", X"00", X"00", X"08", X"00", X"08", X"87", X"77", 
X"9F", X"73", X"F7", X"F9", X"70", X"00", X"08", X"08", X"00", X"00", X"00", X"00", X"08", X"6F", X"76", X"7F", 
X"67", X"76", X"77", X"8F", X"7F", X"FF", X"FF", X"FF", X"FF", X"6F", X"7F", X"FF", X"67", X"27", X"26", X"72", 
X"86", X"27", X"27", X"67", X"72", X"77", X"77", X"67", X"F7", X"77", X"67", X"77", X"7F", X"77", X"88", X"F7", 
X"00", X"68", X"08", X"60", X"86", X"86", X"86", X"86", X"67", X"66", X"76", X"76", X"86", X"06", X"06", X"86", 
X"77", X"C7", X"F6", X"F4", X"F6", X"F6", X"F6", X"F6", X"FC", X"76", X"F6", X"76", X"74", X"00", X"00", X"00", 
X"80", X"00", X"00", X"40", X"40", X"84", X"06", X"06", X"04", X"86", X"06", X"08", X"00", X"00", X"00", X"00", 
X"00", X"08", X"00", X"08", X"06", X"08", X"00", X"00", X"00", X"00", X"00", X"00", X"88", X"88", X"88", X"08", 
X"00", X"80", X"80", X"50", X"88", X"88", X"28", X"73", X"77", X"79", X"79", X"7F", X"78", X"05", X"00", X"04", 
X"00", X"08", X"86", X"86", X"88", X"82", X"67", X"26", X"72", X"67", X"26", X"28", X"37", X"F7", X"F7", X"72", 
X"6E", X"6E", X"7F", X"7F", X"72", X"7E", X"72", X"E7", X"27", X"77", X"E7", X"FE", X"77", X"67", X"77", X"78", 
X"76", X"78", X"77", X"68", X"88", X"77", X"07", X"9F", X"00", X"06", X"80", X"80", X"88", X"62", X"68", X"68", 
X"67", X"67", X"67", X"68", X"68", X"48", X"48", X"67", X"6F", X"77", X"6F", X"67", X"C7", X"66", X"7C", X"76", 
X"6F", X"67", X"C7", X"68", X"80", X"08", X"00", X"60", X"00", X"00", X"00", X"00", X"06", X"08", X"06", X"04", 
X"86", X"86", X"86", X"86", X"00", X"00", X"00", X"80", X"06", X"00", X"06", X"00", X"00", X"08", X"06", X"08", 
X"00", X"08", X"00", X"00", X"88", X"88", X"88", X"00", X"50", X"00", X"00", X"00", X"87", X"88", X"82", X"88", 
X"38", X"73", X"F7", X"79", X"70", X"00", X"00", X"00", X"00", X"00", X"88", X"88", X"26", X"88", X"88", X"28", 
X"78", X"28", X"82", X"87", X"27", X"27", X"27", X"F6", X"27", X"62", X"68", X"82", X"76", X"2F", X"27", X"67", 
X"76", X"27", X"77", X"76", X"72", X"88", X"27", X"23", X"82", X"62", X"82", X"82", X"88", X"83", X"77", X"F7", 
X"08", X"00", X"20", X"68", X"06", X"88", X"67", X"68", X"68", X"67", X"67", X"67", X"68", X"60", X"67", X"7F", 
X"7C", X"7C", X"F6", X"7C", X"F6", X"FC", X"76", X"FC", X"76", X"F6", X"77", X"67", X"40", X"00", X"00", X"00", 
X"08", X"06", X"00", X"80", X"00", X"40", X"40", X"68", X"40", X"60", X"68", X"88", X"00", X"80", X"00", X"00", 
X"00", X"00", X"80", X"06", X"08", X"00", X"00", X"04", X"00", X"04", X"00", X"00", X"88", X"87", X"88", X"00", 
X"00", X"08", X"00", X"88", X"87", X"28", X"88", X"28", X"28", X"28", X"83", X"77", X"78", X"00", X"80", X"08", 
X"00", X"08", X"20", X"20", X"88", X"28", X"28", X"86", X"20", X"68", X"68", X"68", X"88", X"87", X"62", X"77", 
X"62", X"FE", X"62", X"88", X"27", X"76", X"7E", X"72", X"62", X"76", X"26", X"78", X"88", X"28", X"77", X"78", 
X"28", X"88", X"26", X"88", X"28", X"87", X"37", X"F7", X"08", X"00", X"00", X"60", X"80", X"88", X"26", X"86", 
X"86", X"26", X"76", X"86", X"88", X"48", X"7C", X"76", X"7F", X"77", X"CF", X"67", X"C7", X"67", X"C7", X"67", 
X"C7", X"67", X"C7", X"68", X"08", X"00", X"00", X"06", X"00", X"00", X"00", X"00", X"60", X"60", X"40", X"60", 
X"60", X"48", X"86", X"86", X"00", X"00", X"08", X"00", X"80", X"80", X"00", X"08", X"00", X"60", X"88", X"00", 
X"80", X"00", X"08", X"00", X"87", X"57", X"88", X"00", X"80", X"00", X"00", X"88", X"88", X"88", X"87", X"82", 
X"88", X"88", X"08", X"88", X"88", X"80", X"08", X"88", X"80", X"00", X"68", X"60", X"28", X"06", X"08", X"08", 
X"88", X"23", X"82", X"86", X"82", X"87", X"88", X"27", X"76", X"87", X"88", X"28", X"82", X"72", X"72", X"67", 
X"26", X"26", X"23", X"62", X"68", X"82", X"82", X"68", X"28", X"28", X"82", X"86", X"27", X"78", X"F7", X"F7", 
X"80", X"80", X"00", X"80", X"60", X"60", X"67", X"66", X"86", X"76", X"76", X"86", X"86", X"86", X"77", X"F7", 
X"C7", X"6F", X"67", X"C7", X"6F", X"C7", X"6F", X"6F", X"67", X"C7", X"77", X"68", X"06", X"00", X"00", X"00", 
X"00", X"06", X"00", X"40", X"08", X"06", X"04", X"06", X"86", X"86", X"80", X"80", X"00", X"80", X"00", X"00", 
X"00", X"00", X"80", X"00", X"60", X"08", X"00", X"80", X"00", X"80", X"00", X"00", X"87", X"77", X"88", X"00", 
X"05", X"00", X"80", X"88", X"86", X"28", X"88", X"88", X"82", X"88", X"88", X"00", X"00", X"88", X"88", X"67", 
X"88", X"06", X"20", X"28", X"06", X"20", X"28", X"20", X"06", X"88", X"77", X"88", X"88", X"63", X"87", X"88", 
X"28", X"28", X"26", X"82", X"82", X"77", X"6F", X"E6", X"F2", X"F6", X"76", X"88", X"82", X"86", X"77", X"78", 
X"68", X"68", X"28", X"77", X"7F", X"7F", X"7F", X"9F", X"00", X"60", X"80", X"00", X"80", X"88", X"86", X"76", 
X"86", X"86", X"82", X"68", X"68", X"77", X"C7", X"6F", X"6F", X"4F", X"6F", X"6F", X"66", X"F6", X"7C", X"76", 
X"F6", X"76", X"76", X"88", X"00", X"08", X"00", X"06", X"00", X"00", X"00", X"00", X"40", X"40", X"08", X"60", 
X"40", X"68", X"48", X"68", X"00", X"00", X"00", X"80", X"00", X"60", X"08", X"00", X"00", X"06", X"00", X"60", 
X"60", X"00", X"80", X"80", X"87", X"77", X"58", X"80", X"00", X"00", X"00", X"83", X"88", X"88", X"28", X"28", 
X"88", X"28", X"88", X"88", X"80", X"08", X"08", X"82", X"88", X"88", X"80", X"88", X"28", X"88", X"00", X"80", 
X"20", X"82", X"88", X"76", X"78", X"68", X"28", X"28", X"88", X"88", X"88", X"68", X"87", X"72", X"62", X"7E", 
X"6E", X"7E", X"27", X"26", X"80", X"82", X"76", X"28", X"28", X"27", X"67", X"27", X"77", X"F7", X"7F", X"77", 
X"80", X"00", X"00", X"80", X"08", X"00", X"86", X"76", X"86", X"67", X"68", X"86", X"86", X"77", X"F7", X"C7", 
X"6F", X"67", X"C7", X"66", X"F6", X"6F", X"67", X"C7", X"67", X"C7", X"68", X"00", X"60", X"00", X"00", X"00", 
X"00", X"80", X"80", X"80", X"00", X"84", X"60", X"48", X"86", X"88", X"68", X"08", X"00", X"06", X"00", X"00", 
X"80", X"00", X"00", X"60", X"08", X"00", X"08", X"00", X"00", X"60", X"04", X"00", X"79", X"F7", X"88", X"00", 
X"80", X"80", X"08", X"87", X"77", X"82", X"88", X"80", X"28", X"80", X"20", X"88", X"08", X"40", X"08", X"68", 
X"82", X"82", X"82", X"80", X"88", X"20", X"60", X"20", X"86", X"88", X"08", X"88", X"88", X"88", X"88", X"08", 
X"28", X"28", X"28", X"20", X"26", X"37", X"7E", X"67", X"62", X"67", X"E7", X"68", X"82", X"08", X"28", X"26", 
X"78", X"88", X"28", X"7F", X"F7", X"F7", X"F7", X"F7", X"08", X"08", X"00", X"00", X"00", X"60", X"88", X"26", 
X"88", X"68", X"66", X"87", X"F6", X"F6", X"7F", X"6F", X"4F", X"6F", X"6F", X"C7", X"6F", X"4F", X"67", X"7C", 
X"77", X"67", X"76", X"00", X"00", X"00", X"00", X"80", X"00", X"04", X"00", X"00", X"04", X"00", X"06", X"04", 
X"88", X"68", X"86", X"80", X"00", X"00", X"00", X"00", X"00", X"08", X"00", X"06", X"00", X"80", X"60", X"08", 
X"00", X"00", X"00", X"00", X"78", X"78", X"88", X"00", X"00", X"00", X"00", X"87", X"77", X"78", X"67", X"80", 
X"88", X"88", X"80", X"88", X"88", X"88", X"00", X"80", X"80", X"88", X"88", X"62", X"80", X"80", X"00", X"80", 
X"80", X"26", X"28", X"67", X"88", X"26", X"28", X"20", X"88", X"80", X"28", X"88", X"26", X"27", X"62", X"62", 
X"67", X"62", X"67", X"20", X"00", X"08", X"68", X"28", X"62", X"68", X"76", X"77", X"7F", X"7F", X"79", X"F7", 
X"80", X"00", X"06", X"00", X"00", X"00", X"06", X"76", X"86", X"86", X"88", X"67", X"77", X"76", X"F4", X"76", 
X"7C", X"7C", X"76", X"7C", X"7C", X"76", X"C7", X"6F", X"67", X"67", X"40", X"80", X"80", X"00", X"00", X"00", 
X"00", X"00", X"00", X"40", X"00", X"40", X"40", X"06", X"86", X"88", X"40", X"80", X"00", X"00", X"08", X"00", 
X"08", X"00", X"00", X"00", X"06", X"00", X"08", X"06", X"00", X"80", X"08", X"00", X"88", X"78", X"00", X"05", 
X"00", X"80", X"00", X"87", X"77", X"73", X"78", X"28", X"82", X"08", X"78", X"08", X"88", X"28", X"82", X"08", 
X"80", X"28", X"28", X"88", X"26", X"20", X"20", X"80", X"28", X"88", X"08", X"88", X"78", X"88", X"88", X"88", 
X"28", X"68", X"82", X"82", X"08", X"82", X"76", X"76", X"E8", X"68", X"68", X"68", X"60", X"26", X"07", X"60", 
X"68", X"87", X"72", X"F7", X"F7", X"7F", X"7F", X"7F", X"76", X"60", X"00", X"08", X"00", X"80", X"06", X"76", 
X"26", X"06", X"67", X"76", X"7F", X"C7", X"7C", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"76", X"F6", X"7C", 
X"76", X"76", X"80", X"00", X"08", X"00", X"00", X"48", X"00", X"00", X"00", X"08", X"00", X"08", X"06", X"06", 
X"80", X"48", X"80", X"60", X"08", X"00", X"00", X"80", X"00", X"08", X"08", X"00", X"00", X"80", X"60", X"08", 
X"00", X"00", X"40", X"80", X"88", X"81", X"08", X"00", X"00", X"08", X"00", X"87", X"77", X"77", X"77", X"78", 
X"87", X"82", X"82", X"82", X"88", X"68", X"88", X"80", X"00", X"08", X"88", X"28", X"28", X"88", X"02", X"80", 
X"82", X"08", X"02", X"88", X"67", X"78", X"82", X"68", X"02", X"82", X"86", X"82", X"02", X"68", X"72", X"87", 
X"88", X"87", X"76", X"26", X"E6", X"E6", X"26", X"E6", X"67", X"67", X"77", X"F7", X"F7", X"77", X"F9", X"77", 
X"67", X"68", X"80", X"00", X"00", X"08", X"08", X"67", X"68", X"68", X"87", X"7F", X"67", X"76", X"F6", X"7C", 
X"76", X"7C", X"66", X"76", X"6F", X"67", X"C7", X"76", X"76", X"78", X"40", X"00", X"00", X"00", X"00", X"00", 
X"00", X"80", X"08", X"40", X"06", X"04", X"00", X"88", X"48", X"88", X"60", X"80", X"00", X"00", X"00", X"00", 
X"60", X"00", X"00", X"08", X"00", X"00", X"00", X"80", X"06", X"00", X"00", X"80", X"00", X"80", X"80", X"08", 
X"00", X"00", X"08", X"08", X"77", X"77", X"77", X"77", X"88", X"28", X"88", X"88", X"28", X"20", X"08", X"02", 
X"72", X"88", X"26", X"88", X"72", X"72", X"88", X"08", X"80", X"80", X"80", X"82", X"08", X"28", X"88", X"82", 
X"88", X"86", X"88", X"86", X"80", X"82", X"88", X"88", X"88", X"68", X"76", X"E6", X"6E", X"6E", X"6E", X"6E", 
X"7E", X"7F", X"77", X"7F", X"F7", X"79", X"7F", X"7F", X"67", X"66", X"66", X"00", X"80", X"00", X"08", X"76", 
X"86", X"86", X"77", X"C7", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F7", X"CF", X"67", X"C7", X"67", X"67", 
X"47", X"60", X"80", X"60", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"80", X"40", X"48", 
X"88", X"60", X"60", X"80", X"08", X"00", X"00", X"00", X"00", X"00", X"60", X"00", X"80", X"60", X"80", X"60", 
X"00", X"80", X"04", X"08", X"00", X"80", X"80", X"00", X"50", X"80", X"00", X"00", X"87", X"77", X"77", X"77", 
X"78", X"88", X"82", X"68", X"88", X"88", X"28", X"08", X"67", X"20", X"00", X"26", X"82", X"67", X"26", X"28", 
X"28", X"82", X"60", X"80", X"88", X"68", X"28", X"88", X"88", X"87", X"88", X"88", X"88", X"88", X"88", X"68", 
X"88", X"87", X"36", X"7E", X"66", X"F6", X"E6", X"E6", X"E7", X"77", X"7F", X"77", X"78", X"77", X"77", X"7F", 
X"76", X"78", X"88", X"00", X"00", X"00", X"06", X"82", X"68", X"77", X"F6", X"F7", X"C7", X"C7", X"67", X"C7", 
X"C7", X"66", X"C7", X"67", X"6F", X"67", X"C7", X"67", X"76", X"80", X"60", X"00", X"08", X"00", X"00", X"08", 
X"00", X"08", X"00", X"80", X"40", X"04", X"08", X"84", X"84", X"88", X"06", X"00", X"00", X"00", X"00", X"08", 
X"08", X"00", X"00", X"80", X"00", X"08", X"00", X"08", X"00", X"60", X"00", X"00", X"05", X"08", X"80", X"80", 
X"00", X"00", X"80", X"01", X"00", X"88", X"77", X"77", X"77", X"72", X"78", X"77", X"26", X"76", X"86", X"28", 
X"28", X"76", X"28", X"00", X"88", X"28", X"72", X"76", X"78", X"28", X"82", X"08", X"20", X"82", X"08", X"86", 
X"20", X"88", X"67", X"88", X"88", X"88", X"08", X"88", X"77", X"08", X"88", X"66", X"E6", X"E6", X"E6", X"F6", 
X"F7", X"77", X"77", X"77", X"87", X"88", X"88", X"88", X"76", X"66", X"68", X"68", X"00", X"80", X"08", X"67", 
X"76", X"76", X"77", X"76", X"77", X"7C", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"66", X"F6", X"7C", X"76", 
X"76", X"00", X"80", X"00", X"00", X"00", X"00", X"00", X"60", X"00", X"00", X"00", X"00", X"80", X"04", X"08", 
X"88", X"40", X"60", X"80", X"00", X"08", X"00", X"00", X"00", X"80", X"06", X"00", X"60", X"06", X"08", X"06", 
X"00", X"06", X"08", X"08", X"00", X"80", X"50", X"00", X"00", X"10", X"08", X"00", X"80", X"00", X"08", X"88", 
X"77", X"77", X"77", X"77", X"77", X"F7", X"77", X"76", X"72", X"77", X"77", X"28", X"68", X"68", X"68", X"28", 
X"28", X"88", X"86", X"80", X"00", X"08", X"02", X"80", X"86", X"88", X"78", X"86", X"80", X"60", X"00", X"80", 
X"88", X"08", X"68", X"76", X"66", X"E6", X"E6", X"E7", X"E7", X"F7", X"78", X"78", X"78", X"78", X"77", X"F7", 
X"67", X"67", X"68", X"80", X"00", X"00", X"86", X"86", X"77", X"F6", X"FC", X"7C", X"F6", X"76", X"7C", X"76", 
X"6F", X"66", X"66", X"F6", X"F6", X"67", X"67", X"67", X"68", X"00", X"00", X"80", X"00", X"00", X"00", X"00", 
X"00", X"06", X"08", X"40", X"60", X"40", X"88", X"68", X"48", X"88", X"06", X"00", X"08", X"00", X"00", X"80", 
X"00", X"00", X"00", X"00", X"00", X"80", X"00", X"80", X"08", X"00", X"00", X"40", X"08", X"00", X"08", X"08", 
X"00", X"00", X"00", X"00", X"00", X"80", X"00", X"00", X"00", X"88", X"88", X"77", X"77", X"2F", X"7F", X"7F", 
X"F7", X"F7", X"F7", X"F7", X"FF", X"27", X"77", X"77", X"77", X"72", X"77", X"76", X"78", X"76", X"88", X"82", 
X"88", X"88", X"68", X"78", X"80", X"08", X"06", X"08", X"08", X"80", X"86", X"86", X"76", X"6F", X"6F", X"77", 
X"F7", X"77", X"87", X"87", X"88", X"77", X"7F", X"7F", X"76", X"76", X"76", X"86", X"80", X"00", X"08", X"7E", 
X"76", X"77", X"76", X"77", X"CF", X"6F", X"6F", X"C7", X"C7", X"CF", X"7C", X"76", X"76", X"F6", X"76", X"77", 
X"48", X"00", X"60", X"00", X"08", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"04", X"04", X"88", 
X"84", X"84", X"00", X"60", X"00", X"00", X"00", X"06", X"00", X"60", X"80", X"80", X"60", X"08", X"06", X"00", 
X"60", X"06", X"00", X"80", X"08", X"08", X"05", X"00", X"08", X"00", X"80", X"08", X"00", X"08", X"08", X"08", 
X"00", X"00", X"00", X"00", X"88", X"88", X"86", X"86", X"76", X"76", X"76", X"F7", X"77", X"FE", X"FF", X"EF", 
X"FF", X"FF", X"FF", X"FF", X"FF", X"7F", X"FF", X"F7", X"F7", X"F7", X"76", X"F7", X"F6", X"F7", X"77", X"7F", 
X"76", X"F7", X"77", X"77", X"FF", X"7F", X"E7", X"7F", X"78", X"78", X"78", X"88", X"87", X"FF", X"6F", X"7F", 
X"76", X"F7", X"76", X"76", X"80", X"00", X"06", X"77", X"6F", X"6C", X"7F", X"C7", X"67", X"C7", X"76", X"76", 
X"F6", X"76", X"67", X"6F", X"47", X"67", X"67", X"47", X"80", X"00", X"00", X"00", X"00", X"00", X"00", X"80", 
X"00", X"08", X"00", X"60", X"80", X"80", X"80", X"48", X"60", X"80", X"68", X"00", X"00", X"08", X"00", X"00", 
X"00", X"00", X"06", X"00", X"00", X"60", X"00", X"80", X"00", X"80", X"80", X"00", X"00", X"80", X"00", X"80", 
X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"08", X"00", X"00", X"00", X"08", X"08", 
X"08", X"88", X"88", X"86", X"87", X"88", X"88", X"77", X"77", X"77", X"27", X"76", X"F2", X"F6", X"77", X"F7", 
X"E7", X"F7", X"7F", X"6F", X"FF", X"7F", X"FF", X"F7", X"FF", X"FF", X"EF", X"FE", X"7F", X"6F", X"7F", X"F7", 
X"F7", X"77", X"80", X"87", X"7F", X"7F", X"F7", X"F6", X"67", X"76", X"F7", X"76", X"86", X"80", X"87", X"67", 
X"77", X"77", X"67", X"6F", X"6F", X"6F", X"6F", X"66", X"F6", X"6F", X"C7", X"66", X"76", X"7C", X"76", X"86", 
X"80", X"06", X"08", X"00", X"00", X"00", X"00", X"08", X"00", X"04", X"00", X"00", X"04", X"06", X"06", X"08", 
X"48", X"68", X"06", X"00", X"00", X"00", X"00", X"08", X"08", X"00", X"00", X"80", X"80", X"06", X"00", X"68", 
X"06", X"00", X"06", X"88", X"00", X"80", X"80", X"50", X"80", X"05", X"80", X"05", X"08", X"00", X"80", X"08", 
X"00", X"80", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"08", X"08", X"08", X"08", X"88", X"68", X"88", 
X"88", X"86", X"87", X"88", X"88", X"87", X"86", X"88", X"78", X"67", X"67", X"68", X"67", X"67", X"67", X"67", 
X"67", X"67", X"76", X"77", X"77", X"FF", X"7F", X"6F", X"7F", X"FF", X"77", X"7F", X"F7", X"F6", X"F6", X"FF", 
X"7F", X"6F", X"77", X"77", X"67", X"08", X"67", X"77", X"C7", X"CF", X"6F", X"C7", X"67", X"C7", X"C7", X"C7", 
X"C7", X"67", X"6F", X"6F", X"47", X"67", X"67", X"68", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
X"00", X"00", X"08", X"40", X"00", X"00", X"60", X"86", X"88", X"48", X"68", X"00", X"80", X"00", X"80", X"00", 
X"60", X"06", X"00", X"06", X"00", X"80", X"08", X"00", X"00", X"86", X"00", X"04", X"00", X"08", X"00", X"00", 
X"00", X"00", X"00", X"00", X"00", X"05", X"00", X"00", X"00", X"00", X"00", X"80", X"00", X"00", X"00", X"00", 
X"80", X"00", X"00", X"00", X"80", X"00", X"80", X"08", X"88", X"88", X"88", X"88", X"88", X"88", X"88", X"88", 
X"88", X"88", X"88", X"88", X"88", X"88", X"88", X"88", X"80", X"80", X"88", X"7F", X"FF", X"7F", X"6F", X"F7", 
X"F7", X"F7", X"FF", X"7F", X"6F", X"7F", X"7F", X"77", X"77", X"76", X"F6", X"77", X"67", X"68", X"6F", X"67", 
X"77", X"C7", X"67", X"6F", X"6F", X"67", X"6F", X"67", X"6F", X"C7", X"66", X"7C", X"76", X"76", X"77", X"60", 
X"48", X"00", X"00", X"00", X"80", X"00", X"00", X"00", X"80", X"00", X"00", X"08", X"06", X"80", X"48", X"84", 
X"86", X"08", X"06", X"00", X"00", X"00", X"08", X"00", X"00", X"00", X"60", X"00", X"60", X"06", X"00", X"80", 
X"60", X"08", X"08", X"08", X"00", X"80", X"88", X"05", X"08", X"00", X"08", X"00", X"00", X"00", X"08", X"00", 
X"00", X"80", X"00", X"00", X"08", X"00", X"80", X"00", X"00", X"00", X"80", X"00", X"00", X"00", X"08", X"00", 
X"00", X"80", X"80", X"88", X"88", X"80", X"88", X"08", X"00", X"80", X"00", X"00", X"00", X"00", X"00", X"00", 
X"00", X"87", X"7F", X"7F", X"7F", X"7F", X"7F", X"6F", X"7F", X"7F", X"6F", X"7F", X"7F", X"6F", X"6F", X"7F", 
X"7F", X"5F", X"77", X"F6", X"77", X"77", X"67", X"7C", X"76", X"F6", X"FC", X"7C", X"76", X"F6", X"66", X"F6", 
X"67", X"6F", X"67", X"67", X"67", X"C7", X"68", X"80", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
X"00", X"06", X"00", X"40", X"00", X"04", X"08", X"40", X"88", X"48", X"68", X"00", X"08", X"00", X"60", X"00", 
X"80", X"00", X"00", X"80", X"08", X"00", X"60", X"60", X"00", X"80", X"60", X"08", X"00", X"80", X"08", X"00", 
X"00", X"08", X"00", X"08", X"00", X"00", X"00", X"08", X"00", X"00", X"00", X"08", X"00", X"00", X"00", X"00", 
X"00", X"00", X"00", X"00", X"80", X"00", X"00", X"08", X"00", X"00", X"00", X"00", X"00", X"80", X"00", X"80", 
X"08", X"00", X"80", X"00", X"00", X"00", X"00", X"08", X"87", X"7F", X"F7", X"77", X"F6", X"F7", X"F7", X"F7", 
X"F6", X"FF", X"7F", X"6F", X"77", X"F7", X"F7", X"F6", X"C7", X"F4", X"F6", X"77", X"76", X"76", X"F6", X"7F", 
X"67", X"67", X"67", X"77", X"7C", X"6F", X"7C", X"7C", X"F6", X"67", X"C7", X"C7", X"67", X"76", X"76", X"80", 
X"60", X"08", X"00", X"00", X"00", X"08", X"00", X"00", X"00", X"00", X"00", X"00", X"40", X"00", X"80", X"84", 
X"86", X"88", X"86", X"00", X"00", X"00", X"00", X"60", X"00", X"00", X"06", X"08", X"04", X"80", X"00", X"80", 
X"80", X"60", X"06", X"08", X"01", X"08", X"00", X"80", X"80", X"00", X"01", X"00", X"00", X"80", X"00", X"50", 
X"00", X"00", X"80", X"00", X"00", X"00", X"00", X"80", X"08", X"00", X"08", X"00", X"08", X"00", X"80", X"00", 
X"00", X"08", X"00", X"80", X"00", X"08", X"00", X"00", X"00", X"00", X"00", X"80", X"08", X"00", X"88", X"83", 
X"FF", X"77", X"37", X"67", X"FF", X"6F", X"6F", X"6F", X"7F", X"7F", X"7F", X"F6", X"F7", X"7F", X"6F", X"FF", 
X"77", X"77", X"77", X"7C", X"77", X"76", X"7C", X"76", X"FC", X"7C", X"F6", X"C7", X"C7", X"7C", X"67", X"67", 
X"67", X"C7", X"67", X"67", X"67", X"47", X"48", X"00", X"00", X"00", X"00", X"08", X"00", X"00", X"00", X"80", 
X"00", X"00", X"60", X"80", X"80", X"40", X"48", X"08", X"84", X"86", X"88", X"00", X"00", X"00", X"00", X"00", 
X"60", X"08", X"00", X"06", X"00", X"08", X"40", X"04", X"00", X"08", X"08", X"04", X"00", X"80", X"80", X"80", 
X"10", X"00", X"00", X"80", X"80", X"00", X"80", X"00", X"08", X"00", X"00", X"00", X"80", X"08", X"00", X"00", 
X"00", X"08", X"00", X"00", X"00", X"00", X"00", X"80", X"80", X"00", X"00", X"00", X"70", X"00", X"08", X"08", 
X"00", X"08", X"00", X"00", X"00", X"88", X"77", X"FF", X"73", X"78", X"88", X"7F", X"6F", X"F7", X"FF", X"7F", 
X"6F", X"6F", X"F7", X"F7", X"F7", X"FF", X"F7", X"7F", X"FC", X"7F", X"CF", X"77", X"7C", X"7F", X"6F", X"67", 
X"67", X"76", X"F6", X"F6", X"F6", X"6F", X"66", X"F6", X"67", X"67", X"67", X"C7", X"67", X"67", X"80", X"68", 
X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"04", X"00", X"80", X"04", X"04", 
X"88", X"86", X"06", X"06", X"08", X"00", X"80", X"00", X"00", X"00", X"00", X"00", X"06", X"00", X"80", X"80", 
X"60", X"60", X"60", X"08", X"00", X"05", X"08", X"00", X"08", X"08", X"00", X"00", X"05", X"00", X"00", X"00", 
X"00", X"50", X"08", X"00", X"00", X"00", X"00", X"00", X"80", X"00", X"00", X"80", X"08", X"08", X"00", X"00", 
X"00", X"08", X"08", X"07", X"7F", X"77", X"80", X"00", X"80", X"00", X"08", X"08", X"88", X"77", X"7F", X"77", 
X"87", X"87", X"80", X"0F", X"77", X"F6", X"F6", X"F7", X"FF", X"7F", X"7F", X"F6", X"F7", X"F6", X"FF", X"7F", 
X"77", X"77", X"77", X"67", X"67", X"74", X"76", X"F6", X"F6", X"7C", X"76", X"76", X"76", X"F6", X"6F", X"66", 
X"F6", X"76", X"67", X"67", X"C7", X"67", X"68", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
X"80", X"00", X"84", X"00", X"04", X"06", X"06", X"08", X"40", X"86", X"80", X"00", X"00", X"00", X"00", X"80", 
X"00", X"06", X"08", X"06", X"08", X"06", X"06", X"00", X"08", X"00", X"80", X"60", X"88", X"88", X"08", X"80", 
X"80", X"00", X"00", X"00", X"00", X"00", X"80", X"08", X"00", X"00", X"00", X"00", X"80", X"08", X"08", X"00", 
X"00", X"08", X"00", X"00", X"00", X"00", X"50", X"77", X"77", X"77", X"68", X"7F", X"7F", X"7F", X"7F", X"77", 
X"88", X"00", X"80", X"87", X"77", X"FF", X"98", X"87", X"88", X"80", X"08", X"06", X"F6", X"F7", X"FF", X"6F", 
X"6F", X"6F", X"F7", X"FF", X"7F", X"7F", X"7F", X"6F", X"7F", X"C7", X"7C", X"7F", X"C7", X"7C", X"76", X"7C", 
X"76", X"F6", X"76", X"F6", X"67", X"C7", X"66", X"F6", X"67", X"6F", X"67", X"67", X"67", X"86", X"88", X"60", 
X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"08", X"00", X"00", X"80", X"48", 
X"84", X"88", X"60", X"00", X"00", X"60", X"60", X"08", X"00", X"00", X"00", X"00", X"60", X"00", X"08", X"06", 
X"06", X"06", X"08", X"08", X"88", X"87", X"88", X"88", X"88", X"88", X"88", X"88", X"88", X"80", X"88", X"80", 
X"80", X"80", X"05", X"00", X"05", X"00", X"00", X"05", X"00", X"05", X"08", X"00", X"50", X"00", X"08", X"4F", 
X"7F", X"7F", X"7F", X"6F", X"7F", X"6F", X"7F", X"7F", X"7F", X"F7", X"78", X"97", X"F9", X"38", X"77", X"88", 
X"80", X"80", X"00", X"08", X"7F", X"7F", X"6F", X"7F", X"7F", X"F6", X"F7", X"7F", X"7F", X"F7", X"FF", X"7F", 
X"77", X"7F", X"77", X"76", X"76", X"F6", X"FC", X"76", X"F6", X"7C", X"7C", X"76", X"F6", X"76", X"F6", X"67", 
X"F6", X"67", X"67", X"67", X"67", X"68", X"60", X"80", X"08", X"00", X"00", X"00", X"08", X"00", X"00", X"80", 
X"00", X"00", X"00", X"60", X"04", X"04", X"06", X"08", X"48", X"68", X"80", X"00", X"00", X"00", X"00", X"00", 
X"00", X"00", X"84", X"08", X"00", X"60", X"60", X"00", X"00", X"80", X"60", X"06", X"88", X"88", X"87", X"88", 
X"88", X"85", X"88", X"80", X"88", X"88", X"88", X"88", X"88", X"88", X"88", X"88", X"88", X"88", X"88", X"88", 
X"88", X"80", X"80", X"88", X"08", X"08", X"08", X"77", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F6", X"FF", 
X"7F", X"7F", X"F7", X"F7", X"77", X"78", X"88", X"80", X"00", X"00", X"80", X"80", X"76", X"F7", X"F7", X"F6", 
X"F6", X"FF", X"7F", X"F6", X"F7", X"F7", X"F7", X"F7", X"77", X"C7", X"7C", X"77", X"C7", X"67", X"6F", X"67", 
X"C7", X"6F", X"67", X"C6", X"7C", X"7C", X"67", X"C6", X"67", X"67", X"C7", X"67", X"67", X"60", X"60", X"60", 
X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"08", X"00", X"00", X"08", X"00", X"00", X"80", X"60", 
X"88", X"40", X"60", X"00", X"00", X"80", X"00", X"60", X"80", X"00", X"00", X"60", X"80", X"00", X"06", X"06", 
X"06", X"00", X"68", X"08", X"87", X"77", X"87", X"87", X"77", X"78", X"88", X"78", X"88", X"88", X"85", X"88", 
X"85", X"88", X"88", X"88", X"88", X"88", X"88", X"88", X"88", X"88", X"88", X"88", X"88", X"88", X"77", X"76", 
X"77", X"67", X"77", X"F6", X"F7", X"F7", X"F7", X"7F", X"7F", X"77", X"F7", X"FF", X"7F", X"F7", X"F7", X"77", 
X"88", X"00", X"00", X"08", X"8F", X"6F", X"6F", X"7F", X"7F", X"7F", X"67", X"F7", X"FF", X"6F", X"7F", X"7F", 
X"77", X"77", X"C7", X"77", X"76", X"F4", X"76", X"76", X"F6", X"76", X"76", X"F6", X"F6", X"76", X"F6", X"77", 
X"6F", X"67", X"67", X"67", X"76", X"88", X"60", X"60", X"00", X"08", X"00", X"00", X"00", X"80", X"00", X"06", 
X"00", X"00", X"00", X"00", X"40", X"60", X"40", X"60", X"48", X"88", X"40", X"00", X"80", X"00", X"80", X"00", 
X"00", X"00", X"00", X"00", X"60", X"60", X"80", X"08", X"00", X"80", X"00", X"40", X"78", X"87", X"48", X"88", 
X"88", X"88", X"88", X"84", X"88", X"88", X"88", X"88", X"88", X"88", X"88", X"88", X"78", X"48", X"88", X"48", 
X"88", X"78", X"78", X"87", X"87", X"87", X"77", X"77", X"77", X"F7", X"67", X"77", X"76", X"76", X"77", X"67", 
X"76", X"77", X"77", X"77", X"77", X"77", X"77", X"F7", X"77", X"78", X"88", X"08", X"07", X"7F", X"7F", X"6F", 
X"F6", X"FF", X"F7", X"F6", X"F7", X"FF", X"F6", X"F7", X"7C", X"77", X"7C", X"7C", X"7C", X"77", X"C7", X"C7", 
X"67", X"CF", X"67", X"66", X"6F", X"66", X"76", X"67", X"6C", X"76", X"76", X"76", X"76", X"06", X"88", X"06", 
X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"08", 
X"88", X"48", X"80", X"00", X"00", X"60", X"00", X"00", X"00", X"00", X"06", X"80", X"00", X"00", X"60", X"40", 
X"60", X"60", X"68", X"08", X"67", X"77", X"77", X"76", X"77", X"67", X"87", X"87", X"87", X"86", X"88", X"88", 
X"88", X"84", X"88", X"67", X"88", X"88", X"88", X"88", X"68", X"88", X"47", X"88", X"86", X"87", X"6F", X"7F", 
X"7F", X"7F", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F7", X"FF", X"7F", X"7F", X"7F", X"7F", X"77", X"77", 
X"77", X"77", X"77", X"77", X"77", X"76", X"77", X"77", X"77", X"76", X"F6", X"F7", X"F7", X"77", X"F7", X"F7", 
X"77", X"7C", X"77", X"77", X"76", X"F6", X"77", X"76", X"F6", X"66", X"F6", X"F6", X"76", X"6F", X"6F", X"66", 
X"77", X"67", X"C7", X"67", X"68", X"80", X"60", X"60", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
X"80", X"08", X"00", X"08", X"00", X"40", X"04", X"04", X"04", X"08", X"60", X"00", X"60", X"00", X"00", X"00", 
X"80", X"08", X"00", X"06", X"08", X"40", X"00", X"00", X"08", X"06", X"00", X"60", X"FF", X"7F", X"FF", X"7F", 
X"7F", X"7F", X"67", X"77", X"76", X"77", X"76", X"76", X"78", X"78", X"78", X"87", X"78", X"86", X"88", X"78", 
X"88", X"78", X"88", X"76", X"78", X"78", X"87", X"76", X"F6", X"F7", X"76", X"F7", X"F7", X"F7", X"F7", X"F7", 
X"FF", X"7F", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F7", X"F7", X"77", X"77", X"77", X"7F", X"77", X"77", 
X"F6", X"77", X"77", X"76", X"7C", X"F7", X"77", X"77", X"C7", X"77", X"F6", X"7C", X"76", X"7C", X"7C", X"76", 
X"6F", X"76", X"66", X"C7", X"C7", X"66", X"66", X"F6", X"67", X"67", X"67", X"47", X"86", X"80", X"68", X"80", 
X"80", X"00", X"80", X"00", X"08", X"00", X"00", X"00", X"00", X"00", X"00", X"04", X"00", X"80", X"00", X"48", 
X"88", X"68", X"80", X"00", X"08", X"08", X"08", X"00", X"00", X"00", X"00", X"00", X"00", X"08", X"06", X"04", 
X"06", X"00", X"60", X"08", X"66", X"76", X"6F", X"6F", X"6F", X"6F", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", 
X"FF", X"7F", X"7F", X"77", X"F7", X"77", X"77", X"87", X"78", X"78", X"78", X"88", X"88", X"88", X"77", X"77", 
X"77", X"67", X"77", X"77", X"F6", X"F6", X"76", X"F6", X"7F", X"6F", X"67", X"6F", X"67", X"77", X"77", X"77", 
X"F7", X"F7", X"F7", X"F6", X"F7", X"F7", X"FF", X"6F", X"7F", X"FF", X"7F", X"FF", X"F7", X"F6", X"F7", X"F7", 
X"77", X"C7", X"67", X"6F", X"6F", X"67", X"6F", X"67", X"C6", X"6F", X"67", X"76", X"76", X"7C", X"77", X"47", 
X"67", X"C7", X"76", X"76", X"88", X"06", X"08", X"60", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
X"06", X"00", X"00", X"00", X"00", X"04", X"00", X"04", X"86", X"88", X"00", X"00", X"60", X"00", X"00", X"00", 
X"00", X"06", X"06", X"06", X"08", X"60", X"08", X"08", X"00", X"60", X"80", X"60", X"77", X"72", X"77", X"77", 
X"7F", X"67", X"66", X"67", X"67", X"67", X"67", X"67", X"67", X"7F", X"6F", X"FF", X"6F", X"FF", X"FF", X"FF", 
X"FF", X"FF", X"7F", X"F7", X"F7", X"F7", X"77", X"F7", X"77", X"F7", X"F6", X"F6", X"7F", X"7F", X"7F", X"7F", 
X"77", X"F7", X"FF", X"77", X"FF", X"7F", X"7F", X"77", X"77", X"7F", X"6F", X"77", X"F6", X"77", X"77", X"F7", 
X"77", X"76", X"F7", X"77", X"7F", X"7F", X"7F", X"6F", X"77", X"77", X"C7", X"67", X"6F", X"67", X"66", X"F6", 
X"77", X"66", X"F6", X"C7", X"C7", X"67", X"66", X"76", X"76", X"76", X"76", X"76", X"86", X"06", X"08", X"08", 
X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"08", X"00", X"00", X"60", X"00", X"80", X"00", 
X"88", X"46", X"80", X"00", X"00", X"06", X"00", X"80", X"00", X"00", X"00", X"00", X"00", X"80", X"04", X"04", 
X"80", X"60", X"60", X"06", X"27", X"67", X"67", X"62", X"67", X"77", X"77", X"77", X"77", X"77", X"77", X"7F", 
X"67", X"67", X"76", X"67", X"77", X"67", X"6F", X"67", X"6F", X"6F", X"7F", X"FF", X"FF", X"FF", X"FF", X"FF", 
X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"7F", X"7F", X"F7", X"F7", X"7F", X"F7", X"7F", X"67", X"77", X"F6", 
X"F7", X"77", X"77", X"77", X"77", X"F7", X"77", X"77", X"77", X"77", X"67", X"77", X"67", X"76", X"77", X"77", 
X"67", X"C7", X"77", X"C7", X"67", X"CF", X"67", X"C7", X"C6", X"F6", X"67", X"67", X"67", X"67", X"C7", X"6F", 
X"67", X"67", X"67", X"68", X"80", X"00", X"68", X"60", X"00", X"00", X"00", X"00", X"00", X"80", X"00", X"00", 
X"00", X"00", X"00", X"00", X"00", X"04", X"00", X"46", X"04", X"08", X"00", X"08", X"00", X"00", X"00", X"00", 
X"00", X"00", X"08", X"06", X"00", X"06", X"00", X"00", X"60", X"00", X"60", X"80", X"67", X"72", X"77", X"77", 
X"77", X"67", X"76", X"76", X"76", X"76", X"76", X"77", X"77", X"F6", X"77", X"77", X"6F", X"F7", X"77", X"FF", 
X"7F", X"7F", X"6F", X"6F", X"6F", X"6F", X"6F", X"6F", X"7F", X"6F", X"F7", X"F7", X"F6", X"FF", X"FF", X"FC", 
X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F7", X"F7", X"F7", X"7F", X"77", X"77", 
X"77", X"77", X"77", X"77", X"77", X"77", X"77", X"77", X"77", X"7C", X"76", X"F6", X"F6", X"76", X"67", X"67", 
X"67", X"4F", X"66", X"F6", X"7C", X"76", X"76", X"76", X"7C", X"76", X"76", X"86", X"86", X"06", X"08", X"00", 
X"80", X"00", X"00", X"00", X"00", X"00", X"80", X"00", X"00", X"00", X"08", X"00", X"08", X"00", X"00", X"00", 
X"80", X"06", X"00", X"06", X"08", X"00", X"00", X"08", X"00", X"00", X"00", X"00", X"06", X"00", X"06", X"00", 
X"48", X"40", X"06", X"08", X"86", X"76", X"27", X"68", X"27", X"72", X"77", X"77", X"27", X"72", X"77", X"26", 
X"76", X"77", X"76", X"F7", X"76", X"7E", X"76", X"76", X"F6", X"FF", X"6F", X"F7", X"F6", X"FF", X"7F", X"6F", 
X"6F", X"FF", X"6F", X"6F", X"F6", X"F6", X"76", X"7F", X"76", X"6F", X"66", X"F6", X"F7", X"FF", X"7F", X"F7", 
X"FF", X"7F", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", 
X"76", X"77", X"7C", X"76", X"76", X"7C", X"7C", X"76", X"C7", X"66", X"76", X"66", X"76", X"76", X"76", X"76", 
X"76", X"74", X"76", X"86", X"88", X"06", X"06", X"06", X"00", X"00", X"80", X"00", X"00", X"00", X"00", X"08", 
X"00", X"60", X"00", X"00", X"04", X"00", X"40", X"48", X"48", X"06", X"00", X"00", X"00", X"06", X"00", X"00", 
X"00", X"80", X"06", X"00", X"80", X"04", X"80", X"40", X"08", X"06", X"00", X"60", X"72", X"87", X"88", X"88", 
X"86", X"78", X"67", X"67", X"67", X"67", X"67", X"77", X"77", X"76", X"77", X"26", X"77", X"77", X"77", X"7E", 
X"77", X"6F", X"76", X"F6", X"F7", X"67", X"E7", X"F7", X"F6", X"FE", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", 
X"FF", X"FF", X"FF", X"FF", X"E7", X"F6", X"F6", X"F6", X"F6", X"F6", X"76", X"76", X"76", X"76", X"76", X"77", 
X"F6", X"F6", X"F6", X"F6", X"FF", X"6F", X"6F", X"6F", X"F7", X"C7", X"76", X"F4", X"F6", X"76", X"76", X"6F", 
X"67", X"C7", X"C7", X"6F", X"66", X"7C", X"76", X"67", X"67", X"68", X"67", X"06", X"86", X"80", X"60", X"00", 
X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
X"48", X"08", X"00", X"80", X"60", X"00", X"00", X"00", X"00", X"00", X"00", X"60", X"00", X"00", X"60", X"80", 
X"60", X"60", X"80", X"06", X"88", X"27", X"62", X"88", X"88", X"78", X"76", X"77", X"77", X"77", X"67", X"67", 
X"62", X"77", X"67", X"77", X"67", X"67", X"67", X"76", X"77", X"76", X"F7", X"7F", X"6F", X"7F", X"77", X"6F", 
X"67", X"76", X"7E", X"F6", X"FF", X"6F", X"7F", X"FF", X"7F", X"6F", X"6F", X"6F", X"F6", X"FF", X"7F", X"7F", 
X"67", X"77", X"F7", X"77", X"F7", X"77", X"F7", X"67", X"77", X"77", X"77", X"77", X"77", X"67", X"67", X"77", 
X"67", X"76", X"F6", X"76", X"7C", X"76", X"F6", X"76", X"67", X"67", X"67", X"C7", X"67", X"67", X"67", X"7C", 
X"76", X"76", X"78", X"08", X"86", X"82", X"08", X"08", X"00", X"00", X"00", X"08", X"00", X"00", X"80", X"00", 
X"00", X"00", X"04", X"00", X"08", X"08", X"04", X"08", X"00", X"68", X"00", X"40", X"00", X"00", X"80", X"00", 
X"00", X"00", X"00", X"00", X"60", X"80", X"60", X"40", X"40", X"06", X"06", X"00", X"67", X"88", X"88", X"86", 
X"88", X"87", X"88", X"76", X"86", X"78", X"78", X"77", X"78", X"67", X"78", X"67", X"77", X"77", X"76", X"77", 
X"76", X"77", X"67", X"67", X"F7", X"6F", X"6F", X"77", X"F7", X"7F", X"77", X"77", X"7F", X"76", X"F6", X"F6", 
X"F6", X"FF", X"FF", X"7F", X"FF", X"7F", X"F6", X"F7", X"F7", X"6F", X"67", X"76", X"76", X"F6", X"77", X"76", 
X"77", X"67", X"67", X"67", X"77", X"77", X"76", X"77", X"67", X"C7", X"67", X"C7", X"6F", X"66", X"7C", X"7C", 
X"F6", X"7C", X"76", X"76", X"67", X"66", X"76", X"67", X"67", X"68", X"60", X"68", X"00", X"68", X"68", X"06", 
X"08", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"80", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
X"40", X"86", X"00", X"08", X"00", X"00", X"00", X"06", X"00", X"80", X"08", X"00", X"00", X"00", X"68", X"00", 
X"60", X"60", X"00", X"80", X"82", X"86", X"82", X"08", X"82", X"88", X"68", X"87", X"82", X"78", X"62", X"86", 
X"78", X"36", X"78", X"82", X"86", X"82", X"83", X"67", X"27", X"77", X"77", X"F7", X"FF", X"7F", X"7F", X"F6", 
X"F7", X"F6", X"77", X"F6", X"F7", X"FF", X"7F", X"7F", X"7F", X"76", X"F6", X"77", X"6F", X"67", X"77", X"76", 
X"F7", X"77", X"F7", X"77", X"77", X"77", X"67", X"77", X"77", X"77", X"77", X"77", X"67", X"6F", X"77", X"77", 
X"77", X"77", X"C7", X"76", X"67", X"C7", X"66", X"76", X"66", X"76", X"76", X"7C", X"76", X"F6", X"76", X"76", 
X"74", X"76", X"80", X"08", X"80", X"80", X"60", X"80", X"00", X"00", X"80", X"00", X"00", X"00", X"00", X"00", 
X"00", X"08", X"00", X"00", X"04", X"00", X"04", X"08", X"00", X"88", X"00", X"00", X"06", X"00", X"08", X"00", 
X"00", X"04", X"00", X"06", X"06", X"06", X"04", X"06", X"08", X"40", X"60", X"60", X"68", X"82", X"88", X"82", 
X"86", X"87", X"28", X"76", X"87", X"67", X"87", X"87", X"86", X"82", X"82", X"86", X"87", X"87", X"67", X"77", 
X"76", X"27", X"67", X"F7", X"7F", X"7F", X"77", X"F7", X"F6", X"F8", X"FF", X"7F", X"7F", X"6F", X"7F", X"6F", 
X"7F", X"77", X"7F", X"7F", X"77", X"FF", X"7F", X"7F", X"77", X"F7", X"7F", X"6F", X"77", X"7F", X"7F", X"6F", 
X"6F", X"77", X"F6", X"F7", X"F7", X"77", X"6F", X"67", X"4F", X"67", X"76", X"67", X"67", X"66", X"F6", X"76", 
X"76", X"C7", X"66", X"76", X"76", X"67", X"67", X"67", X"68", X"68", X"00", X"06", X"06", X"08", X"06", X"88", 
X"06", X"00", X"00", X"00", X"00", X"80", X"00", X"00", X"00", X"00", X"08", X"00", X"00", X"80", X"00", X"40", 
X"00", X"86", X"80", X"40", X"00", X"00", X"00", X"00", X"00", X"00", X"80", X"00", X"00", X"08", X"04", X"00", 
X"60", X"06", X"00", X"80", X"26", X"77", X"76", X"88", X"82", X"88", X"82", X"88", X"88", X"82", X"86", X"82", 
X"87", X"88", X"78", X"78", X"26", X"78", X"86", X"27", X"77", X"77", X"7E", X"7F", X"6F", X"7F", X"6F", X"7F", 
X"7F", X"77", X"6F", X"6F", X"7F", X"7F", X"7F", X"7F", X"6F", X"77", X"77", X"6F", X"7F", X"6F", X"67", X"77", 
X"F6", X"F6", X"F7", X"F6", X"F6", X"F6", X"77", X"77", X"7F", X"67", X"7F", X"6F", X"7E", X"7F", X"77", X"F7", 
X"76", X"7C", X"76", X"FC", X"76", X"F6", X"66", X"F4", X"76", X"76", X"F6", X"76", X"67", X"67", X"C7", X"67", 
X"68", X"88", X"00", X"88", X"80", X"06", X"00", X"86", X"00", X"00", X"00", X"08", X"00", X"00", X"00", X"00", 
X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"06", X"08", X"60", X"00", X"80", X"00", X"00", X"00", X"00", 
X"00", X"00", X"04", X"00", X"04", X"64", X"80", X"40", X"60", X"60", X"84", X"08", X"88", X"28", X"28", X"87", 
X"88", X"76", X"88", X"72", X"87", X"88", X"82", X"88", X"86", X"86", X"88", X"68", X"78", X"72", X"77", X"86", 
X"76", X"76", X"77", X"77", X"7F", X"7F", X"F7", X"F6", X"F7", X"67", X"F7", X"F7", X"F6", X"F6", X"F7", X"F7", 
X"F7", X"6F", X"77", X"77", X"7F", X"77", X"FF", X"6F", X"7F", X"7F", X"7F", X"7F", X"7F", X"7F", X"F7", X"F6", 
X"F7", X"FF", X"6F", X"77", X"F7", X"76", X"7F", X"67", X"76", X"76", X"76", X"67", X"66", X"7C", X"76", X"67", 
X"C7", X"66", X"76", X"67", X"C7", X"67", X"67", X"47", X"68", X"68", X"00", X"00", X"68", X"00", X"00", X"00", 
X"86", X"00", X"60", X"00", X"00", X"00", X"08", X"00", X"06", X"00", X"00", X"00", X"00", X"00", X"80", X"08", 
X"87", X"84", X"04", X"06", X"04", X"08", X"00", X"00", X"00", X"00", X"00", X"80", X"00", X"06", X"48", X"04", 
X"00", X"40", X"00", X"68", X"88", X"68", X"86", X"82", X"88", X"28", X"78", X"68", X"28", X"67", X"86", X"78", 
X"27", X"87", X"28", X"78", X"87", X"88", X"67", X"72", X"72", X"77", X"7F", X"76", X"7F", X"6F", X"6F", X"7F", 
X"7F", X"8F", X"77", X"6F", X"77", X"77", X"F6", X"F7", X"FF", X"6F", X"6F", X"76", X"F7", X"F6", X"F7", X"F7", 
X"7F", X"7F", X"67", X"6F", X"6F", X"77", X"6F", X"77", X"F6", X"77", X"F7", X"7F", X"6F", X"77", X"F7", X"F7", 
X"7C", X"76", X"7C", X"76", X"7C", X"76", X"7C", X"76", X"67", X"67", X"C7", X"67", X"67", X"67", X"47", X"68", 
X"68", X"00", X"06", X"08", X"00", X"00", X"00", X"80", X"00", X"80", X"00", X"00", X"06", X"00", X"00", X"00", 
X"00", X"00", X"08", X"00", X"00", X"00", X"40", X"04", X"87", X"60", X"80", X"80", X"00", X"00", X"00", X"80", 
X"00", X"08", X"00", X"00", X"48", X"68", X"06", X"08", X"04", X"06", X"08", X"00", X"63", X"82", X"88", X"78", 
X"68", X"88", X"28", X"88", X"88", X"28", X"78", X"28", X"88", X"88", X"88", X"28", X"68", X"72", X"88", X"78", 
X"77", X"76", X"F7", X"7F", X"77", X"7F", X"7F", X"7F", X"77", X"67", X"77", X"7F", X"67", X"F7", X"F7", X"F6", 
X"77", X"77", X"77", X"F7", X"F6", X"F7", X"7F", X"6F", X"6F", X"6F", X"7F", X"77", X"7F", X"6F", X"F6", X"F6", 
X"FF", X"7F", X"6F", X"6F", X"77", X"6F", X"6F", X"77", X"77", X"C7", X"67", X"C6", X"76", X"76", X"76", X"76", 
X"F6", X"67", X"67", X"66", X"74", X"76", X"86", X"86", X"88", X"00", X"00", X"20", X"60", X"80", X"00", X"00", 
X"00", X"08", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"08", X"00", X"00", X"00", X"00", 
X"08", X"04", X"84", X"84", X"80", X"00", X"00", X"08", X"00", X"00", X"80", X"00", X"04", X"86", X"40", X"48", 
X"06", X"08", X"06", X"08", X"88", X"88", X"28", X"28", X"82", X"78", X"86", X"36", X"88", X"82", X"88", X"68", 
X"82", X"63", X"68", X"88", X"28", X"88", X"28", X"28", X"67", X"27", X"F7", X"76", X"77", X"F7", X"F7", X"F6", 
X"F7", X"7F", X"77", X"7F", X"77", X"6F", X"77", X"F7", X"F7", X"77", X"F6", X"77", X"77", X"F7", X"7F", X"77", 
X"7F", X"77", X"7F", X"6F", X"77", X"77", X"77", X"F7", X"7F", X"6F", X"7F", X"77", X"F7", X"77", X"F6", X"F7", 
X"66", X"76", X"76", X"76", X"F6", X"C7", X"C6", X"7C", X"67", X"66", X"76", X"76", X"76", X"76", X"74", X"78", 
X"40", X"08", X"00", X"00", X"00", X"00", X"00", X"60", X"00", X"00", X"06", X"00", X"00", X"00", X"80", X"00", 
X"00", X"80", X"00", X"00", X"00", X"00", X"00", X"40", X"06", X"80", X"60", X"80", X"40", X"00", X"00", X"00", 
X"00", X"00", X"00", X"80", X"86", X"06", X"08", X"04", X"08", X"40", X"00", X"60", X"62", X"78", X"88", X"87", 
X"88", X"68", X"28", X"82", X"86", X"88", X"88", X"78", X"88", X"88", X"87", X"28", X"86", X"78", X"86", X"88", 
X"88", X"77", X"6F", X"77", X"77", X"7F", X"6F", X"7F", X"76", X"7F", X"6F", X"77", X"77", X"F7", X"6F", X"77", 
X"F6", X"F7", X"F7", X"F6", X"F7", X"7C", X"F7", X"7F", X"6F", X"7F", X"67", X"77", X"F6", X"F6", X"F6", X"77", 
X"F6", X"7F", X"77", X"6F", X"6F", X"6F", X"77", X"7F", X"76", X"7C", X"6F", X"66", X"76", X"76", X"F6", X"67", 
X"6F", X"67", X"C7", X"47", X"66", X"86", X"86", X"86", X"08", X"00", X"80", X"88", X"00", X"80", X"00", X"00", 
X"06", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"04", 
X"87", X"68", X"60", X"68", X"04", X"00", X"00", X"00", X"00", X"00", X"04", X"00", X"06", X"86", X"04", X"00", 
X"06", X"06", X"00", X"80", X"88", X"67", X"67", X"62", X"83", X"88", X"88", X"78", X"87", X"82", X"78", X"26", 
X"88", X"28", X"88", X"88", X"88", X"88", X"88", X"78", X"26", X"7F", X"77", X"7F", X"6F", X"7F", X"7F", X"7F", 
X"77", X"77", X"76", X"F7", X"76", X"F7", X"7F", X"67", X"F6", X"7F", X"67", X"7F", X"6F", X"7F", X"6F", X"77", 
X"77", X"6F", X"77", X"76", X"F7", X"F7", X"77", X"67", X"F7", X"6F", X"7F", X"77", X"77", X"7F", X"6F", X"77", 
others => X"00");
end FridgeWelcomeScreen;