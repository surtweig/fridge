(
(X"00", X"00", X"00", X"00", X"00", X"00"), 
(X"7C", X"A2", X"8A", X"A2", X"7C", X"00"), 
(X"7C", X"D6", X"F2", X"D6", X"7C", X"00"), 
(X"38", X"7C", X"3E", X"7C", X"38", X"00"), 
(X"10", X"38", X"7C", X"38", X"10", X"00"), 
(X"18", X"5A", X"FE", X"5A", X"18", X"00"), 
(X"18", X"3A", X"7E", X"3A", X"18", X"00"), 
(X"00", X"18", X"3C", X"3C", X"18", X"00"), 
(X"FF", X"E7", X"C3", X"C3", X"E7", X"FF"), 
(X"00", X"18", X"24", X"24", X"18", X"00"), 
(X"FF", X"E7", X"DB", X"DB", X"E7", X"FF"), 
(X"FE", X"E6", X"CE", X"E6", X"FE", X"00"), 
(X"FE", X"CE", X"E6", X"CE", X"FE", X"00"), 
(X"FE", X"EE", X"C6", X"D6", X"FE", X"00"), 
(X"FE", X"D6", X"C6", X"EE", X"FE", X"00"), 
(X"5A", X"3C", X"E7", X"E7", X"3C", X"5A"), 

(X"7C", X"38", X"38", X"10", X"10", X"00"), 
(X"10", X"10", X"38", X"38", X"7C", X"00"), 
(X"24", X"66", X"FF", X"66", X"24", X"00"), 
(X"00", X"FA", X"00", X"00", X"FA", X"00"), 
(X"60", X"90", X"FE", X"80", X"FE", X"00"), 
(X"5A", X"FD", X"A5", X"BF", X"9A", X"40"), 
(X"00", X"06", X"06", X"06", X"06", X"00"), 
(X"29", X"6D", X"FF", X"FF", X"6D", X"29"), 
(X"20", X"60", X"FE", X"60", X"20", X"00"), 
(X"08", X"0C", X"FE", X"0C", X"08", X"00"), 
(X"10", X"10", X"7C", X"38", X"10", X"00"), 
(X"10", X"38", X"7C", X"10", X"10", X"10"), 
(X"7E", X"46", X"56", X"46", X"7E", X"00"), 
(X"10", X"38", X"10", X"10", X"38", X"10"), 
(X"04", X"1C", X"7C", X"1C", X"04", X"00"), 
(X"40", X"70", X"7C", X"70", X"40", X"00"), 

(X"00", X"00", X"00", X"00", X"00", X"00"), 
(X"00", X"00", X"FA", X"00", X"00", X"00"), 
(X"00", X"20", X"C0", X"20", X"C0", X"00"), 
(X"28", X"FE", X"28", X"FE", X"28", X"00"), 
(X"24", X"54", X"D6", X"54", X"48", X"00"), 
(X"C2", X"0C", X"10", X"60", X"86", X"00"), 
(X"0C", X"52", X"BA", X"4C", X"12", X"00"), 
(X"00", X"00", X"20", X"C0", X"00", X"00"), 
(X"00", X"38", X"44", X"82", X"82", X"00"), 
(X"00", X"82", X"82", X"44", X"38", X"00"), 
(X"00", X"28", X"10", X"10", X"28", X"00"), 
(X"10", X"10", X"7C", X"10", X"10", X"00"), 
(X"00", X"00", X"07", X"00", X"00", X"00"), 
(X"10", X"10", X"10", X"10", X"10", X"00"), 
(X"00", X"00", X"06", X"00", X"00", X"00"), 
(X"02", X"0C", X"10", X"60", X"80", X"00"), 

(X"7C", X"8A", X"92", X"A2", X"7C", X"00"), 
(X"02", X"42", X"FE", X"02", X"02", X"00"), 
(X"46", X"8A", X"92", X"92", X"66", X"00"), 
(X"44", X"82", X"92", X"92", X"6C", X"00"), 
(X"18", X"28", X"48", X"88", X"FE", X"00"), 
(X"E4", X"A2", X"A2", X"A2", X"9C", X"00"), 
(X"3C", X"52", X"92", X"92", X"0C", X"00"), 
(X"C0", X"80", X"8E", X"90", X"E0", X"00"), 
(X"6C", X"92", X"92", X"92", X"6C", X"00"), 
(X"60", X"92", X"92", X"94", X"78", X"00"), 
(X"00", X"00", X"66", X"00", X"00", X"00"), 
(X"00", X"00", X"67", X"00", X"00", X"00"), 
(X"10", X"28", X"44", X"82", X"00", X"00"), 
(X"24", X"24", X"24", X"24", X"24", X"00"), 
(X"82", X"44", X"28", X"10", X"00", X"00"), 
(X"40", X"80", X"8A", X"90", X"60", X"00"), 

(X"7C", X"82", X"BA", X"BA", X"8A", X"78"), 
(X"7E", X"A0", X"A0", X"A0", X"7E", X"00"), 
(X"FE", X"A2", X"A2", X"A2", X"5C", X"00"), 
(X"7C", X"82", X"82", X"82", X"44", X"00"), 
(X"FE", X"82", X"82", X"82", X"7C", X"00"), 
(X"FE", X"A2", X"A2", X"82", X"82", X"00"), 
(X"FE", X"A0", X"A0", X"80", X"80", X"00"), 
(X"7C", X"82", X"82", X"A2", X"BC", X"00"), 
(X"FE", X"20", X"20", X"20", X"FE", X"00"), 
(X"00", X"82", X"FE", X"82", X"00", X"00"), 
(X"04", X"02", X"02", X"02", X"FC", X"00"), 
(X"FE", X"20", X"20", X"50", X"8E", X"00"), 
(X"FE", X"02", X"02", X"02", X"02", X"00"), 
(X"FE", X"40", X"20", X"40", X"FE", X"00"), 
(X"FE", X"40", X"20", X"10", X"FE", X"00"), 
(X"7C", X"82", X"82", X"82", X"7C", X"00"), 

(X"FE", X"A0", X"A0", X"A0", X"40", X"00"), 
(X"7C", X"82", X"82", X"84", X"7A", X"00"), 
(X"FE", X"A0", X"A0", X"A0", X"5E", X"00"), 
(X"44", X"A2", X"A2", X"A2", X"9C", X"00"), 
(X"80", X"80", X"FE", X"80", X"80", X"00"), 
(X"FC", X"02", X"02", X"02", X"FC", X"00"), 
(X"F0", X"0C", X"02", X"0C", X"F0", X"00"), 
(X"FE", X"04", X"08", X"04", X"FE", X"00"), 
(X"8E", X"50", X"20", X"50", X"8E", X"00"), 
(X"80", X"40", X"3E", X"40", X"80", X"00"), 
(X"86", X"8A", X"92", X"A2", X"C2", X"00"), 
(X"00", X"FE", X"82", X"82", X"00", X"00"), 
(X"80", X"60", X"10", X"0C", X"02", X"00"), 
(X"00", X"82", X"82", X"FE", X"00", X"00"), 
(X"20", X"40", X"80", X"40", X"20", X"00"), 
(X"01", X"01", X"01", X"01", X"01", X"00"), 

(X"00", X"00", X"C0", X"20", X"00", X"00"), 
(X"04", X"2A", X"2A", X"2A", X"1E", X"00"), 
(X"FE", X"12", X"22", X"22", X"1C", X"00"), 
(X"1C", X"22", X"22", X"22", X"14", X"00"), 
(X"1C", X"22", X"22", X"12", X"FE", X"00"), 
(X"1C", X"2A", X"2A", X"2A", X"1A", X"00"), 
(X"00", X"20", X"7E", X"A0", X"A0", X"00"), 
(X"19", X"25", X"25", X"25", X"3E", X"00"), 
(X"FE", X"10", X"20", X"20", X"1E", X"00"), 
(X"00", X"00", X"BE", X"00", X"00", X"00"), 
(X"06", X"01", X"01", X"01", X"BE", X"00"), 
(X"00", X"FE", X"08", X"14", X"22", X"00"), 
(X"00", X"00", X"FC", X"02", X"00", X"00"), 
(X"3E", X"20", X"18", X"20", X"1E", X"00"), 
(X"3E", X"20", X"20", X"20", X"1E", X"00"), 
(X"1C", X"22", X"22", X"22", X"1C", X"00"), 

(X"3F", X"14", X"24", X"24", X"18", X"00"), 
(X"18", X"24", X"24", X"14", X"3F", X"00"), 
(X"3E", X"10", X"20", X"20", X"10", X"00"), 
(X"12", X"2A", X"2A", X"2A", X"24", X"00"), 
(X"00", X"20", X"FC", X"22", X"00", X"00"), 
(X"3C", X"02", X"02", X"02", X"3E", X"00"), 
(X"38", X"04", X"02", X"04", X"38", X"00"), 
(X"3C", X"02", X"0E", X"02", X"3E", X"00"), 
(X"22", X"14", X"08", X"14", X"22", X"00"), 
(X"39", X"05", X"05", X"05", X"3E", X"00"), 
(X"22", X"26", X"2A", X"32", X"22", X"00"), 
(X"00", X"10", X"6C", X"82", X"82", X"00"), 
(X"00", X"00", X"EE", X"00", X"00", X"00"), 
(X"00", X"82", X"82", X"6C", X"10", X"00"), 
(X"40", X"80", X"C0", X"40", X"80", X"00"), 
(X"0E", X"12", X"22", X"12", X"0E", X"00"), 

(X"10", X"3E", X"68", X"3E", X"10", X"00"), 
(X"30", X"70", X"7E", X"70", X"30", X"00"), 
(X"44", X"88", X"44", X"11", X"22", X"11"), 
(X"FE", X"FE", X"FE", X"FE", X"FE", X"00"), 
(X"EE", X"EE", X"EE", X"EE", X"EE", X"00"), 
(X"EE", X"EE", X"E0", X"EE", X"EE", X"0E"), 
(X"B5", X"D3", X"CD", X"DE", X"2E", X"B5"), 
(X"FE", X"28", X"EE", X"28", X"FE", X"00"), 
(X"3F", X"F1", X"9F", X"FC", X"C7", X"FF"), 
(X"60", X"06", X"37", X"38", X"83", X"73"), 
(X"FF", X"44", X"44", X"44", X"FF", X"00"), 
(X"44", X"7C", X"44", X"44", X"7C", X"44"), 
(X"0F", X"14", X"24", X"52", X"4B", X"44"), 
(X"4B", X"52", X"24", X"14", X"0F", X"00"), 
(X"E0", X"50", X"48", X"94", X"A4", X"44"), 
(X"A4", X"94", X"48", X"50", X"E0", X"00"), 

(X"FF", X"00", X"18", X"00", X"FF", X"00"), 
(X"44", X"44", X"54", X"54", X"44", X"44"), 
(X"7A", X"58", X"58", X"58", X"7A", X"00"), 
(X"FE", X"BE", X"AA", X"9E", X"FE", X"00"), 
(X"FF", X"88", X"90", X"C2", X"84", X"80"), 
(X"5E", X"5E", X"7E", X"5E", X"5E", X"00"), 
(X"00", X"60", X"9E", X"9E", X"60", X"00"), 
(X"00", X"60", X"FE", X"FE", X"60", X"00"), 
(X"66", X"66", X"16", X"0E", X"06", X"00"), 
(X"06", X"0E", X"16", X"66", X"66", X"00"), 
(X"FE", X"D2", X"92", X"D2", X"FE", X"00"), 
(X"FE", X"AA", X"FE", X"AA", X"FE", X"00"), 
(X"12", X"7E", X"92", X"92", X"42", X"00"), 
(X"7E", X"52", X"66", X"52", X"7E", X"00"), 
(X"00", X"28", X"10", X"28", X"00", X"00"), 
(X"02", X"11", X"7E", X"90", X"40", X"00"), 

(X"7E", X"5E", X"42", X"5E", X"7E", X"00"), 
(X"7E", X"6E", X"42", X"6E", X"7E", X"00"), 
(X"7E", X"76", X"42", X"76", X"7E", X"00"), 
(X"7E", X"7A", X"42", X"7A", X"7E", X"00"), 
(X"22", X"44", X"88", X"44", X"22", X"00"), 
(X"88", X"44", X"22", X"44", X"88", X"00"), 
(X"44", X"28", X"92", X"44", X"28", X"92"), 
(X"92", X"28", X"44", X"92", X"28", X"44"), 
(X"0C", X"12", X"A2", X"02", X"04", X"00"), 
(X"DF", X"9B", X"D9", X"F3", X"BB", X"FE"), 
(X"10", X"10", X"10", X"10", X"1C", X"00"), 
(X"70", X"70", X"76", X"70", X"70", X"00"), 
(X"6E", X"6E", X"66", X"6E", X"6E", X"00"), 
(X"7E", X"72", X"72", X"52", X"7E", X"00"), 
(X"10", X"28", X"54", X"28", X"44", X"00"), 
(X"44", X"28", X"54", X"28", X"10", X"00"), 

(X"AA", X"00", X"55", X"00", X"AA", X"00"), 
(X"AA", X"55", X"AA", X"55", X"AA", X"55"), 
(X"FF", X"55", X"FF", X"AA", X"FF", X"55"), 
(X"00", X"00", X"FF", X"00", X"00", X"00"), 
(X"10", X"10", X"FF", X"00", X"00", X"00"), 
(X"28", X"28", X"FF", X"00", X"00", X"00"), 
(X"10", X"FF", X"00", X"FF", X"00", X"00"), 
(X"10", X"1F", X"10", X"1F", X"00", X"00"), 
(X"28", X"28", X"3F", X"00", X"00", X"00"), 
(X"28", X"EF", X"00", X"FF", X"00", X"00"), 
(X"00", X"FF", X"00", X"FF", X"00", X"00"), 
(X"28", X"2F", X"20", X"3F", X"00", X"00"), 
(X"28", X"E8", X"08", X"F8", X"00", X"00"), 
(X"08", X"F8", X"08", X"F8", X"00", X"00"), 
(X"28", X"28", X"F8", X"00", X"00", X"00"), 
(X"10", X"10", X"1F", X"00", X"00", X"00"), 

(X"00", X"00", X"F0", X"10", X"10", X"10"), 
(X"10", X"10", X"F0", X"10", X"10", X"10"), 
(X"10", X"10", X"1F", X"10", X"10", X"10"), 
(X"00", X"00", X"FF", X"10", X"10", X"10"), 
(X"10", X"10", X"10", X"10", X"10", X"10"), 
(X"10", X"10", X"FF", X"10", X"10", X"10"), 
(X"00", X"00", X"FF", X"28", X"28", X"28"), 
(X"00", X"FF", X"00", X"FF", X"08", X"08"), 
(X"00", X"F8", X"08", X"E8", X"28", X"28"), 
(X"00", X"3F", X"20", X"2F", X"28", X"28"), 
(X"28", X"E8", X"08", X"E8", X"28", X"28"), 
(X"28", X"2F", X"20", X"2F", X"28", X"28"), 
(X"00", X"FF", X"00", X"EF", X"28", X"28"), 
(X"28", X"28", X"28", X"28", X"28", X"28"), 
(X"28", X"EF", X"00", X"EF", X"28", X"28"), 
(X"28", X"28", X"E8", X"28", X"28", X"28"), 

(X"10", X"F0", X"10", X"F0", X"10", X"10"), 
(X"28", X"28", X"2F", X"28", X"28", X"28"), 
(X"10", X"1F", X"10", X"1F", X"10", X"10"), 
(X"00", X"F0", X"10", X"F0", X"10", X"10"), 
(X"00", X"00", X"F8", X"28", X"28", X"28"), 
(X"00", X"00", X"3F", X"28", X"28", X"28"), 
(X"00", X"1F", X"10", X"1F", X"10", X"10"), 
(X"10", X"FF", X"10", X"FF", X"10", X"10"), 
(X"28", X"28", X"FF", X"28", X"28", X"28"), 
(X"10", X"10", X"F0", X"00", X"00", X"00"), 
(X"00", X"00", X"0F", X"08", X"08", X"08"), 
(X"FF", X"FF", X"FF", X"FF", X"FF", X"FF"), 
(X"0F", X"0F", X"0F", X"0F", X"0F", X"0F"), 
(X"FF", X"FF", X"FF", X"00", X"00", X"00"), 
(X"00", X"00", X"00", X"FF", X"FF", X"FF"), 
(X"F0", X"F0", X"F0", X"F0", X"F0", X"F0"), 

(X"FE", X"00", X"FE", X"00", X"FE", X"00"), 
(X"30", X"7E", X"00", X"30", X"7E", X"00"), 
(X"3E", X"2A", X"7A", X"2A", X"3E", X"00"), 
(X"3E", X"3E", X"7E", X"3E", X"3E", X"00"), 
(X"10", X"1E", X"0C", X"0C", X"0E", X"00"), 
(X"18", X"1E", X"1C", X"1C", X"1E", X"00"), 
(X"60", X"7E", X"38", X"38", X"3E", X"00"), 
(X"00", X"10", X"1C", X"0E", X"0C", X"00"), 
(X"76", X"70", X"76", X"70", X"76", X"00"), 
(X"FE", X"92", X"FE", X"92", X"FE", X"00"), 
(X"00", X"00", X"00", X"00", X"00", X"00"), 
(X"00", X"00", X"00", X"00", X"00", X"00"), 
(X"00", X"00", X"00", X"00", X"00", X"00"), 
(X"00", X"00", X"00", X"00", X"00", X"00"), 
(X"00", X"00", X"00", X"00", X"00", X"00"), 
(X"00", X"00", X"00", X"00", X"00", X"00"), 

(X"54", X"54", X"54", X"54", X"54", X"00"), 
(X"22", X"22", X"FA", X"22", X"22", X"00"), 
(X"8A", X"DA", X"72", X"22", X"02", X"00"), 
(X"22", X"72", X"DA", X"8A", X"02", X"00"), 
(X"00", X"00", X"00", X"00", X"00", X"00"), 
(X"00", X"00", X"00", X"00", X"00", X"00"), 
(X"10", X"10", X"54", X"10", X"10", X"00"), 
(X"24", X"48", X"6C", X"24", X"48", X"00"), 
(X"60", X"F0", X"90", X"F0", X"60", X"00"), 
(X"00", X"00", X"18", X"18", X"00", X"00"), 
(X"00", X"00", X"08", X"08", X"00", X"00"), 
(X"08", X"0C", X"06", X"FE", X"80", X"00"), 
(X"F8", X"F8", X"80", X"F8", X"78", X"00"), 
(X"98", X"B8", X"E8", X"48", X"00", X"00"), 
(X"00", X"3C", X"3C", X"3C", X"3C", X"00"), 
(X"00", X"00", X"00", X"00", X"00", X"00")

);